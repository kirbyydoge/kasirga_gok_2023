// Yapay zeka buyruklari
`define MATCH_CNN_LDW   32'h200b
`define MASK_CNN_LDW    32'h7c007fff
`define MATCH_CNN_CLRW  32'h300b
`define MASK_CNN_CLRW   32'hffffffff
`define MATCH_CNN_LDX   32'hb
`define MASK_CNN_LDX    32'h7c007fff
`define MATCH_CNN_CLRX  32'h100b
`define MASK_CNN_CLRX   32'hffffffff
`define MATCH_CNN_RUN   32'h400b
`define MASK_CNN_RUN    32'hfffff07f