`timescale 1ns/1ps

`include "sabitler.vh"
`include "mikroislem.vh"

module dallanma_ongorucu (
     input   [`PS_BIT-1:0]       ps_i,
     input                       ps_gecerli_i,

     output                      ongoru_o, 
     output                      ongoru_gecerli_o


);

endmodule