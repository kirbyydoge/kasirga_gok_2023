`timescale 1ns/1ps

module bellek_islem_birimi(
    input                   clk_i,
    input                   rstn_i
);

endmodule