VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_336x128
   CLASS BLOCK ;
   SIZE 2542.22 BY 583.82 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  556.24 0.0 556.62 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  562.36 0.0 562.74 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  568.48 0.0 568.86 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  573.24 0.0 573.62 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  580.04 0.0 580.42 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  586.16 0.0 586.54 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  591.6 0.0 591.98 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  597.72 0.0 598.1 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  603.84 0.0 604.22 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  609.28 0.0 609.66 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  614.72 0.0 615.1 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  620.84 0.0 621.22 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  626.28 0.0 626.66 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  633.08 0.0 633.46 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  638.52 0.0 638.9 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  644.64 0.0 645.02 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  650.08 0.0 650.46 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  656.2 0.0 656.58 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  661.64 0.0 662.02 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  667.08 0.0 667.46 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  672.52 0.0 672.9 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  678.64 0.0 679.02 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  684.76 0.0 685.14 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  690.2 0.0 690.58 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  696.32 0.0 696.7 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  701.76 0.0 702.14 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  707.88 0.0 708.26 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  714.68 0.0 715.06 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  720.12 0.0 720.5 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  725.56 0.0 725.94 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  732.36 0.0 732.74 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  737.8 0.0 738.18 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  743.24 0.0 743.62 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  748.68 0.0 749.06 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  754.8 0.0 755.18 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  760.92 0.0 761.3 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  767.04 0.0 767.42 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  771.8 0.0 772.18 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  778.6 0.0 778.98 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  784.72 0.0 785.1 1.06 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  790.16 0.0 790.54 1.06 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  796.28 0.0 796.66 1.06 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  801.72 0.0 802.1 1.06 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  807.16 0.0 807.54 1.06 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  813.96 0.0 814.34 1.06 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  818.72 0.0 819.1 1.06 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  825.52 0.0 825.9 1.06 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  830.28 0.0 830.66 1.06 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  837.08 0.0 837.46 1.06 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  843.2 0.0 843.58 1.06 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  848.64 0.0 849.02 1.06 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  854.08 0.0 854.46 1.06 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  860.2 0.0 860.58 1.06 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  866.32 0.0 866.7 1.06 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  872.44 0.0 872.82 1.06 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  877.88 0.0 878.26 1.06 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  883.32 0.0 883.7 1.06 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  889.44 0.0 889.82 1.06 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  894.88 0.0 895.26 1.06 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  901.0 0.0 901.38 1.06 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  907.12 0.0 907.5 1.06 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  912.56 0.0 912.94 1.06 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  918.0 0.0 918.38 1.06 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  924.8 0.0 925.18 1.06 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  929.56 0.0 929.94 1.06 ;
      END
   END din0[64]
   PIN din0[65]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  935.68 0.0 936.06 1.06 ;
      END
   END din0[65]
   PIN din0[66]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  941.8 0.0 942.18 1.06 ;
      END
   END din0[66]
   PIN din0[67]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  947.92 0.0 948.3 1.06 ;
      END
   END din0[67]
   PIN din0[68]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  953.36 0.0 953.74 1.06 ;
      END
   END din0[68]
   PIN din0[69]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  959.48 0.0 959.86 1.06 ;
      END
   END din0[69]
   PIN din0[70]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  965.6 0.0 965.98 1.06 ;
      END
   END din0[70]
   PIN din0[71]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  970.36 0.0 970.74 1.06 ;
      END
   END din0[71]
   PIN din0[72]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  976.48 0.0 976.86 1.06 ;
      END
   END din0[72]
   PIN din0[73]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  983.28 0.0 983.66 1.06 ;
      END
   END din0[73]
   PIN din0[74]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  988.04 0.0 988.42 1.06 ;
      END
   END din0[74]
   PIN din0[75]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  994.84 0.0 995.22 1.06 ;
      END
   END din0[75]
   PIN din0[76]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1000.96 0.0 1001.34 1.06 ;
      END
   END din0[76]
   PIN din0[77]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1006.4 0.0 1006.78 1.06 ;
      END
   END din0[77]
   PIN din0[78]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1011.84 0.0 1012.22 1.06 ;
      END
   END din0[78]
   PIN din0[79]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1017.96 0.0 1018.34 1.06 ;
      END
   END din0[79]
   PIN din0[80]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1023.4 0.0 1023.78 1.06 ;
      END
   END din0[80]
   PIN din0[81]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1030.2 0.0 1030.58 1.06 ;
      END
   END din0[81]
   PIN din0[82]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1035.64 0.0 1036.02 1.06 ;
      END
   END din0[82]
   PIN din0[83]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1041.76 0.0 1042.14 1.06 ;
      END
   END din0[83]
   PIN din0[84]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1047.2 0.0 1047.58 1.06 ;
      END
   END din0[84]
   PIN din0[85]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1053.32 0.0 1053.7 1.06 ;
      END
   END din0[85]
   PIN din0[86]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1058.76 0.0 1059.14 1.06 ;
      END
   END din0[86]
   PIN din0[87]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1064.88 0.0 1065.26 1.06 ;
      END
   END din0[87]
   PIN din0[88]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1071.0 0.0 1071.38 1.06 ;
      END
   END din0[88]
   PIN din0[89]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1076.44 0.0 1076.82 1.06 ;
      END
   END din0[89]
   PIN din0[90]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1081.88 0.0 1082.26 1.06 ;
      END
   END din0[90]
   PIN din0[91]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1088.0 0.0 1088.38 1.06 ;
      END
   END din0[91]
   PIN din0[92]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1094.12 0.0 1094.5 1.06 ;
      END
   END din0[92]
   PIN din0[93]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1098.88 0.0 1099.26 1.06 ;
      END
   END din0[93]
   PIN din0[94]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1105.68 0.0 1106.06 1.06 ;
      END
   END din0[94]
   PIN din0[95]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1111.8 0.0 1112.18 1.06 ;
      END
   END din0[95]
   PIN din0[96]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1116.56 0.0 1116.94 1.06 ;
      END
   END din0[96]
   PIN din0[97]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1123.36 0.0 1123.74 1.06 ;
      END
   END din0[97]
   PIN din0[98]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1128.8 0.0 1129.18 1.06 ;
      END
   END din0[98]
   PIN din0[99]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1134.24 0.0 1134.62 1.06 ;
      END
   END din0[99]
   PIN din0[100]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1140.36 0.0 1140.74 1.06 ;
      END
   END din0[100]
   PIN din0[101]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1146.48 0.0 1146.86 1.06 ;
      END
   END din0[101]
   PIN din0[102]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1152.6 0.0 1152.98 1.06 ;
      END
   END din0[102]
   PIN din0[103]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1158.04 0.0 1158.42 1.06 ;
      END
   END din0[103]
   PIN din0[104]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1163.48 0.0 1163.86 1.06 ;
      END
   END din0[104]
   PIN din0[105]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1169.6 0.0 1169.98 1.06 ;
      END
   END din0[105]
   PIN din0[106]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1175.04 0.0 1175.42 1.06 ;
      END
   END din0[106]
   PIN din0[107]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1181.84 0.0 1182.22 1.06 ;
      END
   END din0[107]
   PIN din0[108]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1187.28 0.0 1187.66 1.06 ;
      END
   END din0[108]
   PIN din0[109]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1193.4 0.0 1193.78 1.06 ;
      END
   END din0[109]
   PIN din0[110]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1198.84 0.0 1199.22 1.06 ;
      END
   END din0[110]
   PIN din0[111]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1204.96 0.0 1205.34 1.06 ;
      END
   END din0[111]
   PIN din0[112]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1211.08 0.0 1211.46 1.06 ;
      END
   END din0[112]
   PIN din0[113]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1216.52 0.0 1216.9 1.06 ;
      END
   END din0[113]
   PIN din0[114]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1222.64 0.0 1223.02 1.06 ;
      END
   END din0[114]
   PIN din0[115]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1227.4 0.0 1227.78 1.06 ;
      END
   END din0[115]
   PIN din0[116]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1234.2 0.0 1234.58 1.06 ;
      END
   END din0[116]
   PIN din0[117]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1239.64 0.0 1240.02 1.06 ;
      END
   END din0[117]
   PIN din0[118]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1245.76 0.0 1246.14 1.06 ;
      END
   END din0[118]
   PIN din0[119]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1251.2 0.0 1251.58 1.06 ;
      END
   END din0[119]
   PIN din0[120]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1257.32 0.0 1257.7 1.06 ;
      END
   END din0[120]
   PIN din0[121]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1263.44 0.0 1263.82 1.06 ;
      END
   END din0[121]
   PIN din0[122]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1268.2 0.0 1268.58 1.06 ;
      END
   END din0[122]
   PIN din0[123]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1275.0 0.0 1275.38 1.06 ;
      END
   END din0[123]
   PIN din0[124]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1281.12 0.0 1281.5 1.06 ;
      END
   END din0[124]
   PIN din0[125]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1286.56 0.0 1286.94 1.06 ;
      END
   END din0[125]
   PIN din0[126]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1292.0 0.0 1292.38 1.06 ;
      END
   END din0[126]
   PIN din0[127]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1298.12 0.0 1298.5 1.06 ;
      END
   END din0[127]
   PIN din0[128]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1303.56 0.0 1303.94 1.06 ;
      END
   END din0[128]
   PIN din0[129]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1309.68 0.0 1310.06 1.06 ;
      END
   END din0[129]
   PIN din0[130]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1315.8 0.0 1316.18 1.06 ;
      END
   END din0[130]
   PIN din0[131]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1321.24 0.0 1321.62 1.06 ;
      END
   END din0[131]
   PIN din0[132]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1328.04 0.0 1328.42 1.06 ;
      END
   END din0[132]
   PIN din0[133]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1332.8 0.0 1333.18 1.06 ;
      END
   END din0[133]
   PIN din0[134]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1339.6 0.0 1339.98 1.06 ;
      END
   END din0[134]
   PIN din0[135]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1345.04 0.0 1345.42 1.06 ;
      END
   END din0[135]
   PIN din0[136]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1351.16 0.0 1351.54 1.06 ;
      END
   END din0[136]
   PIN din0[137]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1355.92 0.0 1356.3 1.06 ;
      END
   END din0[137]
   PIN din0[138]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1362.72 0.0 1363.1 1.06 ;
      END
   END din0[138]
   PIN din0[139]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1368.16 0.0 1368.54 1.06 ;
      END
   END din0[139]
   PIN din0[140]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1373.6 0.0 1373.98 1.06 ;
      END
   END din0[140]
   PIN din0[141]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1379.72 0.0 1380.1 1.06 ;
      END
   END din0[141]
   PIN din0[142]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1385.84 0.0 1386.22 1.06 ;
      END
   END din0[142]
   PIN din0[143]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1391.96 0.0 1392.34 1.06 ;
      END
   END din0[143]
   PIN din0[144]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1398.08 0.0 1398.46 1.06 ;
      END
   END din0[144]
   PIN din0[145]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1403.52 0.0 1403.9 1.06 ;
      END
   END din0[145]
   PIN din0[146]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1409.64 0.0 1410.02 1.06 ;
      END
   END din0[146]
   PIN din0[147]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1415.08 0.0 1415.46 1.06 ;
      END
   END din0[147]
   PIN din0[148]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1421.2 0.0 1421.58 1.06 ;
      END
   END din0[148]
   PIN din0[149]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1427.32 0.0 1427.7 1.06 ;
      END
   END din0[149]
   PIN din0[150]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1432.08 0.0 1432.46 1.06 ;
      END
   END din0[150]
   PIN din0[151]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1438.88 0.0 1439.26 1.06 ;
      END
   END din0[151]
   PIN din0[152]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1444.32 0.0 1444.7 1.06 ;
      END
   END din0[152]
   PIN din0[153]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1450.44 0.0 1450.82 1.06 ;
      END
   END din0[153]
   PIN din0[154]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1455.88 0.0 1456.26 1.06 ;
      END
   END din0[154]
   PIN din0[155]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1462.0 0.0 1462.38 1.06 ;
      END
   END din0[155]
   PIN din0[156]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1468.12 0.0 1468.5 1.06 ;
      END
   END din0[156]
   PIN din0[157]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1473.56 0.0 1473.94 1.06 ;
      END
   END din0[157]
   PIN din0[158]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1479.0 0.0 1479.38 1.06 ;
      END
   END din0[158]
   PIN din0[159]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1484.44 0.0 1484.82 1.06 ;
      END
   END din0[159]
   PIN din0[160]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1491.24 0.0 1491.62 1.06 ;
      END
   END din0[160]
   PIN din0[161]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1496.68 0.0 1497.06 1.06 ;
      END
   END din0[161]
   PIN din0[162]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1502.8 0.0 1503.18 1.06 ;
      END
   END din0[162]
   PIN din0[163]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1508.24 0.0 1508.62 1.06 ;
      END
   END din0[163]
   PIN din0[164]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1514.36 0.0 1514.74 1.06 ;
      END
   END din0[164]
   PIN din0[165]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1519.8 0.0 1520.18 1.06 ;
      END
   END din0[165]
   PIN din0[166]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1525.24 0.0 1525.62 1.06 ;
      END
   END din0[166]
   PIN din0[167]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1531.36 0.0 1531.74 1.06 ;
      END
   END din0[167]
   PIN din0[168]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1537.48 0.0 1537.86 1.06 ;
      END
   END din0[168]
   PIN din0[169]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1542.92 0.0 1543.3 1.06 ;
      END
   END din0[169]
   PIN din0[170]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1549.04 0.0 1549.42 1.06 ;
      END
   END din0[170]
   PIN din0[171]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1554.48 0.0 1554.86 1.06 ;
      END
   END din0[171]
   PIN din0[172]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1560.6 0.0 1560.98 1.06 ;
      END
   END din0[172]
   PIN din0[173]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1566.72 0.0 1567.1 1.06 ;
      END
   END din0[173]
   PIN din0[174]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1572.84 0.0 1573.22 1.06 ;
      END
   END din0[174]
   PIN din0[175]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1578.96 0.0 1579.34 1.06 ;
      END
   END din0[175]
   PIN din0[176]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1583.72 0.0 1584.1 1.06 ;
      END
   END din0[176]
   PIN din0[177]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1590.52 0.0 1590.9 1.06 ;
      END
   END din0[177]
   PIN din0[178]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1595.96 0.0 1596.34 1.06 ;
      END
   END din0[178]
   PIN din0[179]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1601.4 0.0 1601.78 1.06 ;
      END
   END din0[179]
   PIN din0[180]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1608.2 0.0 1608.58 1.06 ;
      END
   END din0[180]
   PIN din0[181]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1612.96 0.0 1613.34 1.06 ;
      END
   END din0[181]
   PIN din0[182]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1619.76 0.0 1620.14 1.06 ;
      END
   END din0[182]
   PIN din0[183]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1625.88 0.0 1626.26 1.06 ;
      END
   END din0[183]
   PIN din0[184]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1631.32 0.0 1631.7 1.06 ;
      END
   END din0[184]
   PIN din0[185]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1636.76 0.0 1637.14 1.06 ;
      END
   END din0[185]
   PIN din0[186]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1642.88 0.0 1643.26 1.06 ;
      END
   END din0[186]
   PIN din0[187]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1648.32 0.0 1648.7 1.06 ;
      END
   END din0[187]
   PIN din0[188]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1654.44 0.0 1654.82 1.06 ;
      END
   END din0[188]
   PIN din0[189]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1660.56 0.0 1660.94 1.06 ;
      END
   END din0[189]
   PIN din0[190]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1665.32 0.0 1665.7 1.06 ;
      END
   END din0[190]
   PIN din0[191]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1672.12 0.0 1672.5 1.06 ;
      END
   END din0[191]
   PIN din0[192]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1677.56 0.0 1677.94 1.06 ;
      END
   END din0[192]
   PIN din0[193]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1683.68 0.0 1684.06 1.06 ;
      END
   END din0[193]
   PIN din0[194]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1689.8 0.0 1690.18 1.06 ;
      END
   END din0[194]
   PIN din0[195]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1695.24 0.0 1695.62 1.06 ;
      END
   END din0[195]
   PIN din0[196]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1701.36 0.0 1701.74 1.06 ;
      END
   END din0[196]
   PIN din0[197]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1706.8 0.0 1707.18 1.06 ;
      END
   END din0[197]
   PIN din0[198]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1712.92 0.0 1713.3 1.06 ;
      END
   END din0[198]
   PIN din0[199]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1719.04 0.0 1719.42 1.06 ;
      END
   END din0[199]
   PIN din0[200]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1725.16 0.0 1725.54 1.06 ;
      END
   END din0[200]
   PIN din0[201]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1730.6 0.0 1730.98 1.06 ;
      END
   END din0[201]
   PIN din0[202]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1736.72 0.0 1737.1 1.06 ;
      END
   END din0[202]
   PIN din0[203]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1741.48 0.0 1741.86 1.06 ;
      END
   END din0[203]
   PIN din0[204]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1748.28 0.0 1748.66 1.06 ;
      END
   END din0[204]
   PIN din0[205]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1753.04 0.0 1753.42 1.06 ;
      END
   END din0[205]
   PIN din0[206]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1759.84 0.0 1760.22 1.06 ;
      END
   END din0[206]
   PIN din0[207]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1765.28 0.0 1765.66 1.06 ;
      END
   END din0[207]
   PIN din0[208]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1771.4 0.0 1771.78 1.06 ;
      END
   END din0[208]
   PIN din0[209]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1776.84 0.0 1777.22 1.06 ;
      END
   END din0[209]
   PIN din0[210]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1782.96 0.0 1783.34 1.06 ;
      END
   END din0[210]
   PIN din0[211]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1788.4 0.0 1788.78 1.06 ;
      END
   END din0[211]
   PIN din0[212]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1795.2 0.0 1795.58 1.06 ;
      END
   END din0[212]
   PIN din0[213]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1799.96 0.0 1800.34 1.06 ;
      END
   END din0[213]
   PIN din0[214]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1806.08 0.0 1806.46 1.06 ;
      END
   END din0[214]
   PIN din0[215]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1812.2 0.0 1812.58 1.06 ;
      END
   END din0[215]
   PIN din0[216]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1817.64 0.0 1818.02 1.06 ;
      END
   END din0[216]
   PIN din0[217]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1823.08 0.0 1823.46 1.06 ;
      END
   END din0[217]
   PIN din0[218]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1829.88 0.0 1830.26 1.06 ;
      END
   END din0[218]
   PIN din0[219]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1836.0 0.0 1836.38 1.06 ;
      END
   END din0[219]
   PIN din0[220]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1841.44 0.0 1841.82 1.06 ;
      END
   END din0[220]
   PIN din0[221]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1846.88 0.0 1847.26 1.06 ;
      END
   END din0[221]
   PIN din0[222]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1853.0 0.0 1853.38 1.06 ;
      END
   END din0[222]
   PIN din0[223]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1859.12 0.0 1859.5 1.06 ;
      END
   END din0[223]
   PIN din0[224]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1863.88 0.0 1864.26 1.06 ;
      END
   END din0[224]
   PIN din0[225]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1870.68 0.0 1871.06 1.06 ;
      END
   END din0[225]
   PIN din0[226]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1876.8 0.0 1877.18 1.06 ;
      END
   END din0[226]
   PIN din0[227]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1881.56 0.0 1881.94 1.06 ;
      END
   END din0[227]
   PIN din0[228]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1888.36 0.0 1888.74 1.06 ;
      END
   END din0[228]
   PIN din0[229]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1893.12 0.0 1893.5 1.06 ;
      END
   END din0[229]
   PIN din0[230]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1899.92 0.0 1900.3 1.06 ;
      END
   END din0[230]
   PIN din0[231]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1906.04 0.0 1906.42 1.06 ;
      END
   END din0[231]
   PIN din0[232]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1911.48 0.0 1911.86 1.06 ;
      END
   END din0[232]
   PIN din0[233]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1916.92 0.0 1917.3 1.06 ;
      END
   END din0[233]
   PIN din0[234]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1922.36 0.0 1922.74 1.06 ;
      END
   END din0[234]
   PIN din0[235]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1928.48 0.0 1928.86 1.06 ;
      END
   END din0[235]
   PIN din0[236]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1934.6 0.0 1934.98 1.06 ;
      END
   END din0[236]
   PIN din0[237]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1940.04 0.0 1940.42 1.06 ;
      END
   END din0[237]
   PIN din0[238]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1946.16 0.0 1946.54 1.06 ;
      END
   END din0[238]
   PIN din0[239]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1951.6 0.0 1951.98 1.06 ;
      END
   END din0[239]
   PIN din0[240]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1957.72 0.0 1958.1 1.06 ;
      END
   END din0[240]
   PIN din0[241]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1963.16 0.0 1963.54 1.06 ;
      END
   END din0[241]
   PIN din0[242]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1969.28 0.0 1969.66 1.06 ;
      END
   END din0[242]
   PIN din0[243]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1976.08 0.0 1976.46 1.06 ;
      END
   END din0[243]
   PIN din0[244]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1980.84 0.0 1981.22 1.06 ;
      END
   END din0[244]
   PIN din0[245]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1986.96 0.0 1987.34 1.06 ;
      END
   END din0[245]
   PIN din0[246]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1993.08 0.0 1993.46 1.06 ;
      END
   END din0[246]
   PIN din0[247]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1998.52 0.0 1998.9 1.06 ;
      END
   END din0[247]
   PIN din0[248]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2004.64 0.0 2005.02 1.06 ;
      END
   END din0[248]
   PIN din0[249]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2010.76 0.0 2011.14 1.06 ;
      END
   END din0[249]
   PIN din0[250]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2016.88 0.0 2017.26 1.06 ;
      END
   END din0[250]
   PIN din0[251]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2023.0 0.0 2023.38 1.06 ;
      END
   END din0[251]
   PIN din0[252]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2028.44 0.0 2028.82 1.06 ;
      END
   END din0[252]
   PIN din0[253]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2034.56 0.0 2034.94 1.06 ;
      END
   END din0[253]
   PIN din0[254]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2040.0 0.0 2040.38 1.06 ;
      END
   END din0[254]
   PIN din0[255]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2046.12 0.0 2046.5 1.06 ;
      END
   END din0[255]
   PIN din0[256]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2050.88 0.0 2051.26 1.06 ;
      END
   END din0[256]
   PIN din0[257]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2057.68 0.0 2058.06 1.06 ;
      END
   END din0[257]
   PIN din0[258]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2062.44 0.0 2062.82 1.06 ;
      END
   END din0[258]
   PIN din0[259]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2069.24 0.0 2069.62 1.06 ;
      END
   END din0[259]
   PIN din0[260]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2074.68 0.0 2075.06 1.06 ;
      END
   END din0[260]
   PIN din0[261]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2080.8 0.0 2081.18 1.06 ;
      END
   END din0[261]
   PIN din0[262]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2086.24 0.0 2086.62 1.06 ;
      END
   END din0[262]
   PIN din0[263]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2092.36 0.0 2092.74 1.06 ;
      END
   END din0[263]
   PIN din0[264]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2097.8 0.0 2098.18 1.06 ;
      END
   END din0[264]
   PIN din0[265]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2103.92 0.0 2104.3 1.06 ;
      END
   END din0[265]
   PIN din0[266]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2109.36 0.0 2109.74 1.06 ;
      END
   END din0[266]
   PIN din0[267]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2116.16 0.0 2116.54 1.06 ;
      END
   END din0[267]
   PIN din0[268]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2122.28 0.0 2122.66 1.06 ;
      END
   END din0[268]
   PIN din0[269]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2127.72 0.0 2128.1 1.06 ;
      END
   END din0[269]
   PIN din0[270]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2133.16 0.0 2133.54 1.06 ;
      END
   END din0[270]
   PIN din0[271]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2139.28 0.0 2139.66 1.06 ;
      END
   END din0[271]
   PIN din0[272]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2144.72 0.0 2145.1 1.06 ;
      END
   END din0[272]
   PIN din0[273]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2150.84 0.0 2151.22 1.06 ;
      END
   END din0[273]
   PIN din0[274]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2156.28 0.0 2156.66 1.06 ;
      END
   END din0[274]
   PIN din0[275]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2162.4 0.0 2162.78 1.06 ;
      END
   END din0[275]
   PIN din0[276]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2167.84 0.0 2168.22 1.06 ;
      END
   END din0[276]
   PIN din0[277]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2173.96 0.0 2174.34 1.06 ;
      END
   END din0[277]
   PIN din0[278]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2180.08 0.0 2180.46 1.06 ;
      END
   END din0[278]
   PIN din0[279]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2185.52 0.0 2185.9 1.06 ;
      END
   END din0[279]
   PIN din0[280]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2191.64 0.0 2192.02 1.06 ;
      END
   END din0[280]
   PIN din0[281]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2197.08 0.0 2197.46 1.06 ;
      END
   END din0[281]
   PIN din0[282]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2203.88 0.0 2204.26 1.06 ;
      END
   END din0[282]
   PIN din0[283]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2208.64 0.0 2209.02 1.06 ;
      END
   END din0[283]
   PIN din0[284]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2214.76 0.0 2215.14 1.06 ;
      END
   END din0[284]
   PIN din0[285]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2220.2 0.0 2220.58 1.06 ;
      END
   END din0[285]
   PIN din0[286]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2226.32 0.0 2226.7 1.06 ;
      END
   END din0[286]
   PIN din0[287]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2233.12 0.0 2233.5 1.06 ;
      END
   END din0[287]
   PIN din0[288]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2237.88 0.0 2238.26 1.06 ;
      END
   END din0[288]
   PIN din0[289]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2244.68 0.0 2245.06 1.06 ;
      END
   END din0[289]
   PIN din0[290]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2249.44 0.0 2249.82 1.06 ;
      END
   END din0[290]
   PIN din0[291]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2256.24 0.0 2256.62 1.06 ;
      END
   END din0[291]
   PIN din0[292]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2261.0 0.0 2261.38 1.06 ;
      END
   END din0[292]
   PIN din0[293]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2267.8 0.0 2268.18 1.06 ;
      END
   END din0[293]
   PIN din0[294]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2273.24 0.0 2273.62 1.06 ;
      END
   END din0[294]
   PIN din0[295]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2279.36 0.0 2279.74 1.06 ;
      END
   END din0[295]
   PIN din0[296]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2285.48 0.0 2285.86 1.06 ;
      END
   END din0[296]
   PIN din0[297]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2290.92 0.0 2291.3 1.06 ;
      END
   END din0[297]
   PIN din0[298]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2297.04 0.0 2297.42 1.06 ;
      END
   END din0[298]
   PIN din0[299]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2303.16 0.0 2303.54 1.06 ;
      END
   END din0[299]
   PIN din0[300]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2308.6 0.0 2308.98 1.06 ;
      END
   END din0[300]
   PIN din0[301]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2314.72 0.0 2315.1 1.06 ;
      END
   END din0[301]
   PIN din0[302]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2320.16 0.0 2320.54 1.06 ;
      END
   END din0[302]
   PIN din0[303]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2326.28 0.0 2326.66 1.06 ;
      END
   END din0[303]
   PIN din0[304]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2331.72 0.0 2332.1 1.06 ;
      END
   END din0[304]
   PIN din0[305]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2337.84 0.0 2338.22 1.06 ;
      END
   END din0[305]
   PIN din0[306]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2343.96 0.0 2344.34 1.06 ;
      END
   END din0[306]
   PIN din0[307]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2348.72 0.0 2349.1 1.06 ;
      END
   END din0[307]
   PIN din0[308]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2355.52 0.0 2355.9 1.06 ;
      END
   END din0[308]
   PIN din0[309]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2360.28 0.0 2360.66 1.06 ;
      END
   END din0[309]
   PIN din0[310]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2366.4 0.0 2366.78 1.06 ;
      END
   END din0[310]
   PIN din0[311]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2372.52 0.0 2372.9 1.06 ;
      END
   END din0[311]
   PIN din0[312]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2377.96 0.0 2378.34 1.06 ;
      END
   END din0[312]
   PIN din0[313]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2384.76 0.0 2385.14 1.06 ;
      END
   END din0[313]
   PIN din0[314]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2390.88 0.0 2391.26 1.06 ;
      END
   END din0[314]
   PIN din0[315]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2396.32 0.0 2396.7 1.06 ;
      END
   END din0[315]
   PIN din0[316]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2401.76 0.0 2402.14 1.06 ;
      END
   END din0[316]
   PIN din0[317]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2407.88 0.0 2408.26 1.06 ;
      END
   END din0[317]
   PIN din0[318]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2413.32 0.0 2413.7 1.06 ;
      END
   END din0[318]
   PIN din0[319]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2418.76 0.0 2419.14 1.06 ;
      END
   END din0[319]
   PIN din0[320]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2424.88 0.0 2425.26 1.06 ;
      END
   END din0[320]
   PIN din0[321]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2431.0 0.0 2431.38 1.06 ;
      END
   END din0[321]
   PIN din0[322]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2437.12 0.0 2437.5 1.06 ;
      END
   END din0[322]
   PIN din0[323]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2442.56 0.0 2442.94 1.06 ;
      END
   END din0[323]
   PIN din0[324]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2448.0 0.0 2448.38 1.06 ;
      END
   END din0[324]
   PIN din0[325]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2454.8 0.0 2455.18 1.06 ;
      END
   END din0[325]
   PIN din0[326]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2460.92 0.0 2461.3 1.06 ;
      END
   END din0[326]
   PIN din0[327]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2466.36 0.0 2466.74 1.06 ;
      END
   END din0[327]
   PIN din0[328]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2471.8 0.0 2472.18 1.06 ;
      END
   END din0[328]
   PIN din0[329]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2477.92 0.0 2478.3 1.06 ;
      END
   END din0[329]
   PIN din0[330]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2483.36 0.0 2483.74 1.06 ;
      END
   END din0[330]
   PIN din0[331]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2489.48 0.0 2489.86 1.06 ;
      END
   END din0[331]
   PIN din0[332]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2494.92 0.0 2495.3 1.06 ;
      END
   END din0[332]
   PIN din0[333]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2501.72 0.0 2502.1 1.06 ;
      END
   END din0[333]
   PIN din0[334]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2506.48 0.0 2506.86 1.06 ;
      END
   END din0[334]
   PIN din0[335]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2513.28 0.0 2513.66 1.06 ;
      END
   END din0[335]
   PIN din0[336]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2519.4 0.0 2519.78 1.06 ;
      END
   END din0[336]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 582.76 296.86 583.82 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 582.76 302.98 583.82 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.16 582.76 297.54 583.82 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.92 582.76 302.3 583.82 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 582.76 301.62 583.82 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 582.76 298.22 583.82 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 582.76 300.94 583.82 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  299.88 582.76 300.26 583.82 ;
      END
   END addr0[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 280.16 1.06 280.54 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 288.32 1.06 288.7 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 280.84 1.06 281.22 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 0.0 311.82 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  316.88 0.0 317.26 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 0.0 323.38 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  328.44 0.0 328.82 1.06 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  334.56 0.0 334.94 1.06 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  340.0 0.0 340.38 1.06 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  346.8 0.0 347.18 1.06 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  351.56 0.0 351.94 1.06 ;
      END
   END wmask0[7]
   PIN wmask0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  358.36 0.0 358.74 1.06 ;
      END
   END wmask0[8]
   PIN wmask0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  363.12 0.0 363.5 1.06 ;
      END
   END wmask0[9]
   PIN wmask0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  369.92 0.0 370.3 1.06 ;
      END
   END wmask0[10]
   PIN wmask0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  376.04 0.0 376.42 1.06 ;
      END
   END wmask0[11]
   PIN wmask0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  381.48 0.0 381.86 1.06 ;
      END
   END wmask0[12]
   PIN wmask0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  386.92 0.0 387.3 1.06 ;
      END
   END wmask0[13]
   PIN wmask0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  393.04 0.0 393.42 1.06 ;
      END
   END wmask0[14]
   PIN wmask0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  398.48 0.0 398.86 1.06 ;
      END
   END wmask0[15]
   PIN wmask0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  405.28 0.0 405.66 1.06 ;
      END
   END wmask0[16]
   PIN wmask0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  410.04 0.0 410.42 1.06 ;
      END
   END wmask0[17]
   PIN wmask0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  416.84 0.0 417.22 1.06 ;
      END
   END wmask0[18]
   PIN wmask0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  421.6 0.0 421.98 1.06 ;
      END
   END wmask0[19]
   PIN wmask0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  428.4 0.0 428.78 1.06 ;
      END
   END wmask0[20]
   PIN wmask0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  433.16 0.0 433.54 1.06 ;
      END
   END wmask0[21]
   PIN wmask0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  439.96 0.0 440.34 1.06 ;
      END
   END wmask0[22]
   PIN wmask0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  445.4 0.0 445.78 1.06 ;
      END
   END wmask0[23]
   PIN wmask0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  451.52 0.0 451.9 1.06 ;
      END
   END wmask0[24]
   PIN wmask0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  456.96 0.0 457.34 1.06 ;
      END
   END wmask0[25]
   PIN wmask0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  463.08 0.0 463.46 1.06 ;
      END
   END wmask0[26]
   PIN wmask0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  469.2 0.0 469.58 1.06 ;
      END
   END wmask0[27]
   PIN wmask0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  475.32 0.0 475.7 1.06 ;
      END
   END wmask0[28]
   PIN wmask0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  480.76 0.0 481.14 1.06 ;
      END
   END wmask0[29]
   PIN wmask0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  486.88 0.0 487.26 1.06 ;
      END
   END wmask0[30]
   PIN wmask0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  491.64 0.0 492.02 1.06 ;
      END
   END wmask0[31]
   PIN wmask0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  498.44 0.0 498.82 1.06 ;
      END
   END wmask0[32]
   PIN wmask0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  503.2 0.0 503.58 1.06 ;
      END
   END wmask0[33]
   PIN wmask0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  510.0 0.0 510.38 1.06 ;
      END
   END wmask0[34]
   PIN wmask0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  515.44 0.0 515.82 1.06 ;
      END
   END wmask0[35]
   PIN wmask0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  520.88 0.0 521.26 1.06 ;
      END
   END wmask0[36]
   PIN wmask0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  527.68 0.0 528.06 1.06 ;
      END
   END wmask0[37]
   PIN wmask0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  533.8 0.0 534.18 1.06 ;
      END
   END wmask0[38]
   PIN wmask0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  539.24 0.0 539.62 1.06 ;
      END
   END wmask0[39]
   PIN wmask0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  544.68 0.0 545.06 1.06 ;
      END
   END wmask0[40]
   PIN wmask0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  550.12 0.0 550.5 1.06 ;
      END
   END wmask0[41]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  2524.84 0.0 2525.22 1.06 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  378.08 582.76 378.46 583.82 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  382.16 582.76 382.54 583.82 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  383.52 582.76 383.9 583.82 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  386.24 582.76 386.62 583.82 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  388.28 582.76 388.66 583.82 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  391.68 582.76 392.06 583.82 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  393.72 582.76 394.1 583.82 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  396.44 582.76 396.82 583.82 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  397.8 582.76 398.18 583.82 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  402.56 582.76 402.94 583.82 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  403.24 582.76 403.62 583.82 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  407.32 582.76 407.7 583.82 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  408.0 582.76 408.38 583.82 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  411.4 582.76 411.78 583.82 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 582.76 413.14 583.82 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 582.76 417.9 583.82 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  418.88 582.76 419.26 583.82 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  422.28 582.76 422.66 583.82 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  422.96 582.76 423.34 583.82 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  426.36 582.76 426.74 583.82 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  427.72 582.76 428.1 583.82 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  432.48 582.76 432.86 583.82 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  433.84 582.76 434.22 583.82 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  436.56 582.76 436.94 583.82 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  437.92 582.76 438.3 583.82 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.0 582.76 442.38 583.82 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  443.36 582.76 443.74 583.82 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  447.44 582.76 447.82 583.82 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  448.12 582.76 448.5 583.82 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  451.52 582.76 451.9 583.82 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  452.88 582.76 453.26 583.82 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  456.28 582.76 456.66 583.82 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  457.64 582.76 458.02 583.82 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  462.4 582.76 462.78 583.82 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  463.08 582.76 463.46 583.82 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.16 582.76 467.54 583.82 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  467.84 582.76 468.22 583.82 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  471.24 582.76 471.62 583.82 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  472.6 582.76 472.98 583.82 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  477.36 582.76 477.74 583.82 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  478.72 582.76 479.1 583.82 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  482.12 582.76 482.5 583.82 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  483.48 582.76 483.86 583.82 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  487.56 582.76 487.94 583.82 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  488.24 582.76 488.62 583.82 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  491.64 582.76 492.02 583.82 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  493.68 582.76 494.06 583.82 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  496.4 582.76 496.78 583.82 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  497.76 582.76 498.14 583.82 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  501.84 582.76 502.22 583.82 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  503.2 582.76 503.58 583.82 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  507.28 582.76 507.66 583.82 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  507.96 582.76 508.34 583.82 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  511.36 582.76 511.74 583.82 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  513.4 582.76 513.78 583.82 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  517.48 582.76 517.86 583.82 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  518.84 582.76 519.22 583.82 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  521.56 582.76 521.94 583.82 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  522.92 582.76 523.3 583.82 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  526.32 582.76 526.7 583.82 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  527.68 582.76 528.06 583.82 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  531.76 582.76 532.14 583.82 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  533.12 582.76 533.5 583.82 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  536.52 582.76 536.9 583.82 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  538.56 582.76 538.94 583.82 ;
      END
   END dout0[64]
   PIN dout0[65]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  541.28 582.76 541.66 583.82 ;
      END
   END dout0[65]
   PIN dout0[66]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  542.64 582.76 543.02 583.82 ;
      END
   END dout0[66]
   PIN dout0[67]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  547.4 582.76 547.78 583.82 ;
      END
   END dout0[67]
   PIN dout0[68]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  548.08 582.76 548.46 583.82 ;
      END
   END dout0[68]
   PIN dout0[69]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  551.48 582.76 551.86 583.82 ;
      END
   END dout0[69]
   PIN dout0[70]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  552.84 582.76 553.22 583.82 ;
      END
   END dout0[70]
   PIN dout0[71]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  556.24 582.76 556.62 583.82 ;
      END
   END dout0[71]
   PIN dout0[72]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  557.6 582.76 557.98 583.82 ;
      END
   END dout0[72]
   PIN dout0[73]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  561.68 582.76 562.06 583.82 ;
      END
   END dout0[73]
   PIN dout0[74]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  563.04 582.76 563.42 583.82 ;
      END
   END dout0[74]
   PIN dout0[75]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  566.44 582.76 566.82 583.82 ;
      END
   END dout0[75]
   PIN dout0[76]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  567.8 582.76 568.18 583.82 ;
      END
   END dout0[76]
   PIN dout0[77]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  572.56 582.76 572.94 583.82 ;
      END
   END dout0[77]
   PIN dout0[78]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  573.24 582.76 573.62 583.82 ;
      END
   END dout0[78]
   PIN dout0[79]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  577.32 582.76 577.7 583.82 ;
      END
   END dout0[79]
   PIN dout0[80]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  578.68 582.76 579.06 583.82 ;
      END
   END dout0[80]
   PIN dout0[81]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  581.4 582.76 581.78 583.82 ;
      END
   END dout0[81]
   PIN dout0[82]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  582.76 582.76 583.14 583.82 ;
      END
   END dout0[82]
   PIN dout0[83]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  587.52 582.76 587.9 583.82 ;
      END
   END dout0[83]
   PIN dout0[84]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  588.2 582.76 588.58 583.82 ;
      END
   END dout0[84]
   PIN dout0[85]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  591.6 582.76 591.98 583.82 ;
      END
   END dout0[85]
   PIN dout0[86]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  592.96 582.76 593.34 583.82 ;
      END
   END dout0[86]
   PIN dout0[87]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  596.36 582.76 596.74 583.82 ;
      END
   END dout0[87]
   PIN dout0[88]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  598.4 582.76 598.78 583.82 ;
      END
   END dout0[88]
   PIN dout0[89]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  602.48 582.76 602.86 583.82 ;
      END
   END dout0[89]
   PIN dout0[90]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  603.16 582.76 603.54 583.82 ;
      END
   END dout0[90]
   PIN dout0[91]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  607.24 582.76 607.62 583.82 ;
      END
   END dout0[91]
   PIN dout0[92]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  607.92 582.76 608.3 583.82 ;
      END
   END dout0[92]
   PIN dout0[93]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  611.32 582.76 611.7 583.82 ;
      END
   END dout0[93]
   PIN dout0[94]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 582.76 613.06 583.82 ;
      END
   END dout0[94]
   PIN dout0[95]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  617.44 582.76 617.82 583.82 ;
      END
   END dout0[95]
   PIN dout0[96]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  618.8 582.76 619.18 583.82 ;
      END
   END dout0[96]
   PIN dout0[97]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  622.2 582.76 622.58 583.82 ;
      END
   END dout0[97]
   PIN dout0[98]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  623.56 582.76 623.94 583.82 ;
      END
   END dout0[98]
   PIN dout0[99]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  626.96 582.76 627.34 583.82 ;
      END
   END dout0[99]
   PIN dout0[100]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  627.64 582.76 628.02 583.82 ;
      END
   END dout0[100]
   PIN dout0[101]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  631.72 582.76 632.1 583.82 ;
      END
   END dout0[101]
   PIN dout0[102]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  633.08 582.76 633.46 583.82 ;
      END
   END dout0[102]
   PIN dout0[103]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  636.48 582.76 636.86 583.82 ;
      END
   END dout0[103]
   PIN dout0[104]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  638.52 582.76 638.9 583.82 ;
      END
   END dout0[104]
   PIN dout0[105]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  641.24 582.76 641.62 583.82 ;
      END
   END dout0[105]
   PIN dout0[106]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  643.28 582.76 643.66 583.82 ;
      END
   END dout0[106]
   PIN dout0[107]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  646.68 582.76 647.06 583.82 ;
      END
   END dout0[107]
   PIN dout0[108]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  648.04 582.76 648.42 583.82 ;
      END
   END dout0[108]
   PIN dout0[109]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  651.44 582.76 651.82 583.82 ;
      END
   END dout0[109]
   PIN dout0[110]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  652.8 582.76 653.18 583.82 ;
      END
   END dout0[110]
   PIN dout0[111]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  657.56 582.76 657.94 583.82 ;
      END
   END dout0[111]
   PIN dout0[112]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  658.24 582.76 658.62 583.82 ;
      END
   END dout0[112]
   PIN dout0[113]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  662.32 582.76 662.7 583.82 ;
      END
   END dout0[113]
   PIN dout0[114]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  663.68 582.76 664.06 583.82 ;
      END
   END dout0[114]
   PIN dout0[115]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  667.08 582.76 667.46 583.82 ;
      END
   END dout0[115]
   PIN dout0[116]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  667.76 582.76 668.14 583.82 ;
      END
   END dout0[116]
   PIN dout0[117]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  672.52 582.76 672.9 583.82 ;
      END
   END dout0[117]
   PIN dout0[118]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  673.88 582.76 674.26 583.82 ;
      END
   END dout0[118]
   PIN dout0[119]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  677.28 582.76 677.66 583.82 ;
      END
   END dout0[119]
   PIN dout0[120]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  678.64 582.76 679.02 583.82 ;
      END
   END dout0[120]
   PIN dout0[121]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  681.36 582.76 681.74 583.82 ;
      END
   END dout0[121]
   PIN dout0[122]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  682.72 582.76 683.1 583.82 ;
      END
   END dout0[122]
   PIN dout0[123]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  686.8 582.76 687.18 583.82 ;
      END
   END dout0[123]
   PIN dout0[124]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  688.16 582.76 688.54 583.82 ;
      END
   END dout0[124]
   PIN dout0[125]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  691.56 582.76 691.94 583.82 ;
      END
   END dout0[125]
   PIN dout0[126]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  692.92 582.76 693.3 583.82 ;
      END
   END dout0[126]
   PIN dout0[127]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  697.0 582.76 697.38 583.82 ;
      END
   END dout0[127]
   PIN dout0[128]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  698.36 582.76 698.74 583.82 ;
      END
   END dout0[128]
   PIN dout0[129]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  702.44 582.76 702.82 583.82 ;
      END
   END dout0[129]
   PIN dout0[130]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  703.12 582.76 703.5 583.82 ;
      END
   END dout0[130]
   PIN dout0[131]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  706.52 582.76 706.9 583.82 ;
      END
   END dout0[131]
   PIN dout0[132]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  707.88 582.76 708.26 583.82 ;
      END
   END dout0[132]
   PIN dout0[133]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  711.28 582.76 711.66 583.82 ;
      END
   END dout0[133]
   PIN dout0[134]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  712.64 582.76 713.02 583.82 ;
      END
   END dout0[134]
   PIN dout0[135]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  717.4 582.76 717.78 583.82 ;
      END
   END dout0[135]
   PIN dout0[136]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  718.08 582.76 718.46 583.82 ;
      END
   END dout0[136]
   PIN dout0[137]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  721.48 582.76 721.86 583.82 ;
      END
   END dout0[137]
   PIN dout0[138]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  722.84 582.76 723.22 583.82 ;
      END
   END dout0[138]
   PIN dout0[139]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  726.24 582.76 726.62 583.82 ;
      END
   END dout0[139]
   PIN dout0[140]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  728.28 582.76 728.66 583.82 ;
      END
   END dout0[140]
   PIN dout0[141]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  732.36 582.76 732.74 583.82 ;
      END
   END dout0[141]
   PIN dout0[142]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  733.04 582.76 733.42 583.82 ;
      END
   END dout0[142]
   PIN dout0[143]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  736.44 582.76 736.82 583.82 ;
      END
   END dout0[143]
   PIN dout0[144]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  737.8 582.76 738.18 583.82 ;
      END
   END dout0[144]
   PIN dout0[145]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  742.56 582.76 742.94 583.82 ;
      END
   END dout0[145]
   PIN dout0[146]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  743.24 582.76 743.62 583.82 ;
      END
   END dout0[146]
   PIN dout0[147]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  746.64 582.76 747.02 583.82 ;
      END
   END dout0[147]
   PIN dout0[148]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  748.0 582.76 748.38 583.82 ;
      END
   END dout0[148]
   PIN dout0[149]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  752.08 582.76 752.46 583.82 ;
      END
   END dout0[149]
   PIN dout0[150]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  752.76 582.76 753.14 583.82 ;
      END
   END dout0[150]
   PIN dout0[151]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  756.84 582.76 757.22 583.82 ;
      END
   END dout0[151]
   PIN dout0[152]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  758.88 582.76 759.26 583.82 ;
      END
   END dout0[152]
   PIN dout0[153]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  762.28 582.76 762.66 583.82 ;
      END
   END dout0[153]
   PIN dout0[154]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  762.96 582.76 763.34 583.82 ;
      END
   END dout0[154]
   PIN dout0[155]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  766.36 582.76 766.74 583.82 ;
      END
   END dout0[155]
   PIN dout0[156]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  767.72 582.76 768.1 583.82 ;
      END
   END dout0[156]
   PIN dout0[157]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  771.8 582.76 772.18 583.82 ;
      END
   END dout0[157]
   PIN dout0[158]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  773.16 582.76 773.54 583.82 ;
      END
   END dout0[158]
   PIN dout0[159]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  776.56 582.76 776.94 583.82 ;
      END
   END dout0[159]
   PIN dout0[160]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  777.92 582.76 778.3 583.82 ;
      END
   END dout0[160]
   PIN dout0[161]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  782.0 582.76 782.38 583.82 ;
      END
   END dout0[161]
   PIN dout0[162]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  782.68 582.76 783.06 583.82 ;
      END
   END dout0[162]
   PIN dout0[163]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  786.76 582.76 787.14 583.82 ;
      END
   END dout0[163]
   PIN dout0[164]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  788.12 582.76 788.5 583.82 ;
      END
   END dout0[164]
   PIN dout0[165]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  791.52 582.76 791.9 583.82 ;
      END
   END dout0[165]
   PIN dout0[166]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  792.88 582.76 793.26 583.82 ;
      END
   END dout0[166]
   PIN dout0[167]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  796.28 582.76 796.66 583.82 ;
      END
   END dout0[167]
   PIN dout0[168]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  797.64 582.76 798.02 583.82 ;
      END
   END dout0[168]
   PIN dout0[169]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  802.4 582.76 802.78 583.82 ;
      END
   END dout0[169]
   PIN dout0[170]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  803.08 582.76 803.46 583.82 ;
      END
   END dout0[170]
   PIN dout0[171]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  806.48 582.76 806.86 583.82 ;
      END
   END dout0[171]
   PIN dout0[172]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  807.84 582.76 808.22 583.82 ;
      END
   END dout0[172]
   PIN dout0[173]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  811.24 582.76 811.62 583.82 ;
      END
   END dout0[173]
   PIN dout0[174]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  813.28 582.76 813.66 583.82 ;
      END
   END dout0[174]
   PIN dout0[175]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  816.68 582.76 817.06 583.82 ;
      END
   END dout0[175]
   PIN dout0[176]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  818.72 582.76 819.1 583.82 ;
      END
   END dout0[176]
   PIN dout0[177]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  822.12 582.76 822.5 583.82 ;
      END
   END dout0[177]
   PIN dout0[178]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  822.8 582.76 823.18 583.82 ;
      END
   END dout0[178]
   PIN dout0[179]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  827.56 582.76 827.94 583.82 ;
      END
   END dout0[179]
   PIN dout0[180]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  828.24 582.76 828.62 583.82 ;
      END
   END dout0[180]
   PIN dout0[181]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  831.64 582.76 832.02 583.82 ;
      END
   END dout0[181]
   PIN dout0[182]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  833.0 582.76 833.38 583.82 ;
      END
   END dout0[182]
   PIN dout0[183]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  836.4 582.76 836.78 583.82 ;
      END
   END dout0[183]
   PIN dout0[184]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  837.76 582.76 838.14 583.82 ;
      END
   END dout0[184]
   PIN dout0[185]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  842.52 582.76 842.9 583.82 ;
      END
   END dout0[185]
   PIN dout0[186]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  843.2 582.76 843.58 583.82 ;
      END
   END dout0[186]
   PIN dout0[187]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  846.6 582.76 846.98 583.82 ;
      END
   END dout0[187]
   PIN dout0[188]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  847.96 582.76 848.34 583.82 ;
      END
   END dout0[188]
   PIN dout0[189]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  851.36 582.76 851.74 583.82 ;
      END
   END dout0[189]
   PIN dout0[190]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  852.72 582.76 853.1 583.82 ;
      END
   END dout0[190]
   PIN dout0[191]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  857.48 582.76 857.86 583.82 ;
      END
   END dout0[191]
   PIN dout0[192]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  858.84 582.76 859.22 583.82 ;
      END
   END dout0[192]
   PIN dout0[193]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  862.24 582.76 862.62 583.82 ;
      END
   END dout0[193]
   PIN dout0[194]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  862.92 582.76 863.3 583.82 ;
      END
   END dout0[194]
   PIN dout0[195]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  866.32 582.76 866.7 583.82 ;
      END
   END dout0[195]
   PIN dout0[196]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  867.68 582.76 868.06 583.82 ;
      END
   END dout0[196]
   PIN dout0[197]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  871.76 582.76 872.14 583.82 ;
      END
   END dout0[197]
   PIN dout0[198]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  873.12 582.76 873.5 583.82 ;
      END
   END dout0[198]
   PIN dout0[199]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  877.2 582.76 877.58 583.82 ;
      END
   END dout0[199]
   PIN dout0[200]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  877.88 582.76 878.26 583.82 ;
      END
   END dout0[200]
   PIN dout0[201]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  881.28 582.76 881.66 583.82 ;
      END
   END dout0[201]
   PIN dout0[202]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  883.32 582.76 883.7 583.82 ;
      END
   END dout0[202]
   PIN dout0[203]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  887.4 582.76 887.78 583.82 ;
      END
   END dout0[203]
   PIN dout0[204]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  888.08 582.76 888.46 583.82 ;
      END
   END dout0[204]
   PIN dout0[205]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  891.48 582.76 891.86 583.82 ;
      END
   END dout0[205]
   PIN dout0[206]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  892.84 582.76 893.22 583.82 ;
      END
   END dout0[206]
   PIN dout0[207]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  896.24 582.76 896.62 583.82 ;
      END
   END dout0[207]
   PIN dout0[208]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  898.28 582.76 898.66 583.82 ;
      END
   END dout0[208]
   PIN dout0[209]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  901.68 582.76 902.06 583.82 ;
      END
   END dout0[209]
   PIN dout0[210]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  903.04 582.76 903.42 583.82 ;
      END
   END dout0[210]
   PIN dout0[211]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  906.44 582.76 906.82 583.82 ;
      END
   END dout0[211]
   PIN dout0[212]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  907.8 582.76 908.18 583.82 ;
      END
   END dout0[212]
   PIN dout0[213]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  911.88 582.76 912.26 583.82 ;
      END
   END dout0[213]
   PIN dout0[214]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  913.24 582.76 913.62 583.82 ;
      END
   END dout0[214]
   PIN dout0[215]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  916.64 582.76 917.02 583.82 ;
      END
   END dout0[215]
   PIN dout0[216]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  918.0 582.76 918.38 583.82 ;
      END
   END dout0[216]
   PIN dout0[217]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  921.4 582.76 921.78 583.82 ;
      END
   END dout0[217]
   PIN dout0[218]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  923.44 582.76 923.82 583.82 ;
      END
   END dout0[218]
   PIN dout0[219]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  927.52 582.76 927.9 583.82 ;
      END
   END dout0[219]
   PIN dout0[220]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  928.2 582.76 928.58 583.82 ;
      END
   END dout0[220]
   PIN dout0[221]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  931.6 582.76 931.98 583.82 ;
      END
   END dout0[221]
   PIN dout0[222]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  932.96 582.76 933.34 583.82 ;
      END
   END dout0[222]
   PIN dout0[223]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  936.36 582.76 936.74 583.82 ;
      END
   END dout0[223]
   PIN dout0[224]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  937.72 582.76 938.1 583.82 ;
      END
   END dout0[224]
   PIN dout0[225]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  941.8 582.76 942.18 583.82 ;
      END
   END dout0[225]
   PIN dout0[226]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  943.16 582.76 943.54 583.82 ;
      END
   END dout0[226]
   PIN dout0[227]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  947.24 582.76 947.62 583.82 ;
      END
   END dout0[227]
   PIN dout0[228]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  947.92 582.76 948.3 583.82 ;
      END
   END dout0[228]
   PIN dout0[229]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  952.0 582.76 952.38 583.82 ;
      END
   END dout0[229]
   PIN dout0[230]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  952.68 582.76 953.06 583.82 ;
      END
   END dout0[230]
   PIN dout0[231]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  957.44 582.76 957.82 583.82 ;
      END
   END dout0[231]
   PIN dout0[232]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  958.8 582.76 959.18 583.82 ;
      END
   END dout0[232]
   PIN dout0[233]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  961.52 582.76 961.9 583.82 ;
      END
   END dout0[233]
   PIN dout0[234]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  963.56 582.76 963.94 583.82 ;
      END
   END dout0[234]
   PIN dout0[235]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  966.96 582.76 967.34 583.82 ;
      END
   END dout0[235]
   PIN dout0[236]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  968.32 582.76 968.7 583.82 ;
      END
   END dout0[236]
   PIN dout0[237]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  971.72 582.76 972.1 583.82 ;
      END
   END dout0[237]
   PIN dout0[238]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  973.08 582.76 973.46 583.82 ;
      END
   END dout0[238]
   PIN dout0[239]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  976.48 582.76 976.86 583.82 ;
      END
   END dout0[239]
   PIN dout0[240]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  977.84 582.76 978.22 583.82 ;
      END
   END dout0[240]
   PIN dout0[241]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  981.92 582.76 982.3 583.82 ;
      END
   END dout0[241]
   PIN dout0[242]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  983.28 582.76 983.66 583.82 ;
      END
   END dout0[242]
   PIN dout0[243]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  986.68 582.76 987.06 583.82 ;
      END
   END dout0[243]
   PIN dout0[244]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  988.04 582.76 988.42 583.82 ;
      END
   END dout0[244]
   PIN dout0[245]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  991.44 582.76 991.82 583.82 ;
      END
   END dout0[245]
   PIN dout0[246]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  992.8 582.76 993.18 583.82 ;
      END
   END dout0[246]
   PIN dout0[247]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  997.56 582.76 997.94 583.82 ;
      END
   END dout0[247]
   PIN dout0[248]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  998.24 582.76 998.62 583.82 ;
      END
   END dout0[248]
   PIN dout0[249]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1001.64 582.76 1002.02 583.82 ;
      END
   END dout0[249]
   PIN dout0[250]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1003.0 582.76 1003.38 583.82 ;
      END
   END dout0[250]
   PIN dout0[251]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1007.08 582.76 1007.46 583.82 ;
      END
   END dout0[251]
   PIN dout0[252]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1008.44 582.76 1008.82 583.82 ;
      END
   END dout0[252]
   PIN dout0[253]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1012.52 582.76 1012.9 583.82 ;
      END
   END dout0[253]
   PIN dout0[254]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1013.88 582.76 1014.26 583.82 ;
      END
   END dout0[254]
   PIN dout0[255]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1016.6 582.76 1016.98 583.82 ;
      END
   END dout0[255]
   PIN dout0[256]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1017.96 582.76 1018.34 583.82 ;
      END
   END dout0[256]
   PIN dout0[257]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1021.36 582.76 1021.74 583.82 ;
      END
   END dout0[257]
   PIN dout0[258]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1022.72 582.76 1023.1 583.82 ;
      END
   END dout0[258]
   PIN dout0[259]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1027.48 582.76 1027.86 583.82 ;
      END
   END dout0[259]
   PIN dout0[260]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1028.16 582.76 1028.54 583.82 ;
      END
   END dout0[260]
   PIN dout0[261]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1032.24 582.76 1032.62 583.82 ;
      END
   END dout0[261]
   PIN dout0[262]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1032.92 582.76 1033.3 583.82 ;
      END
   END dout0[262]
   PIN dout0[263]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1037.0 582.76 1037.38 583.82 ;
      END
   END dout0[263]
   PIN dout0[264]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1038.36 582.76 1038.74 583.82 ;
      END
   END dout0[264]
   PIN dout0[265]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1041.76 582.76 1042.14 583.82 ;
      END
   END dout0[265]
   PIN dout0[266]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1043.8 582.76 1044.18 583.82 ;
      END
   END dout0[266]
   PIN dout0[267]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1047.2 582.76 1047.58 583.82 ;
      END
   END dout0[267]
   PIN dout0[268]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1047.88 582.76 1048.26 583.82 ;
      END
   END dout0[268]
   PIN dout0[269]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1051.28 582.76 1051.66 583.82 ;
      END
   END dout0[269]
   PIN dout0[270]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1053.32 582.76 1053.7 583.82 ;
      END
   END dout0[270]
   PIN dout0[271]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1057.4 582.76 1057.78 583.82 ;
      END
   END dout0[271]
   PIN dout0[272]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1058.08 582.76 1058.46 583.82 ;
      END
   END dout0[272]
   PIN dout0[273]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1061.48 582.76 1061.86 583.82 ;
      END
   END dout0[273]
   PIN dout0[274]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1062.84 582.76 1063.22 583.82 ;
      END
   END dout0[274]
   PIN dout0[275]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1066.92 582.76 1067.3 583.82 ;
      END
   END dout0[275]
   PIN dout0[276]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1068.28 582.76 1068.66 583.82 ;
      END
   END dout0[276]
   PIN dout0[277]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1071.68 582.76 1072.06 583.82 ;
      END
   END dout0[277]
   PIN dout0[278]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1073.04 582.76 1073.42 583.82 ;
      END
   END dout0[278]
   PIN dout0[279]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1076.44 582.76 1076.82 583.82 ;
      END
   END dout0[279]
   PIN dout0[280]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1078.48 582.76 1078.86 583.82 ;
      END
   END dout0[280]
   PIN dout0[281]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1082.56 582.76 1082.94 583.82 ;
      END
   END dout0[281]
   PIN dout0[282]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1083.92 582.76 1084.3 583.82 ;
      END
   END dout0[282]
   PIN dout0[283]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1087.32 582.76 1087.7 583.82 ;
      END
   END dout0[283]
   PIN dout0[284]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1088.0 582.76 1088.38 583.82 ;
      END
   END dout0[284]
   PIN dout0[285]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1091.4 582.76 1091.78 583.82 ;
      END
   END dout0[285]
   PIN dout0[286]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1092.76 582.76 1093.14 583.82 ;
      END
   END dout0[286]
   PIN dout0[287]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1097.52 582.76 1097.9 583.82 ;
      END
   END dout0[287]
   PIN dout0[288]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1098.2 582.76 1098.58 583.82 ;
      END
   END dout0[288]
   PIN dout0[289]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1102.28 582.76 1102.66 583.82 ;
      END
   END dout0[289]
   PIN dout0[290]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1103.64 582.76 1104.02 583.82 ;
      END
   END dout0[290]
   PIN dout0[291]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1107.04 582.76 1107.42 583.82 ;
      END
   END dout0[291]
   PIN dout0[292]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1108.4 582.76 1108.78 583.82 ;
      END
   END dout0[292]
   PIN dout0[293]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1112.48 582.76 1112.86 583.82 ;
      END
   END dout0[293]
   PIN dout0[294]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1113.16 582.76 1113.54 583.82 ;
      END
   END dout0[294]
   PIN dout0[295]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1116.56 582.76 1116.94 583.82 ;
      END
   END dout0[295]
   PIN dout0[296]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1118.6 582.76 1118.98 583.82 ;
      END
   END dout0[296]
   PIN dout0[297]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1121.32 582.76 1121.7 583.82 ;
      END
   END dout0[297]
   PIN dout0[298]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1122.68 582.76 1123.06 583.82 ;
      END
   END dout0[298]
   PIN dout0[299]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1126.76 582.76 1127.14 583.82 ;
      END
   END dout0[299]
   PIN dout0[300]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1128.12 582.76 1128.5 583.82 ;
      END
   END dout0[300]
   PIN dout0[301]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1131.52 582.76 1131.9 583.82 ;
      END
   END dout0[301]
   PIN dout0[302]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1132.88 582.76 1133.26 583.82 ;
      END
   END dout0[302]
   PIN dout0[303]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1136.28 582.76 1136.66 583.82 ;
      END
   END dout0[303]
   PIN dout0[304]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1138.32 582.76 1138.7 583.82 ;
      END
   END dout0[304]
   PIN dout0[305]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1142.4 582.76 1142.78 583.82 ;
      END
   END dout0[305]
   PIN dout0[306]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1143.76 582.76 1144.14 583.82 ;
      END
   END dout0[306]
   PIN dout0[307]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1146.48 582.76 1146.86 583.82 ;
      END
   END dout0[307]
   PIN dout0[308]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1147.84 582.76 1148.22 583.82 ;
      END
   END dout0[308]
   PIN dout0[309]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1151.24 582.76 1151.62 583.82 ;
      END
   END dout0[309]
   PIN dout0[310]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1152.6 582.76 1152.98 583.82 ;
      END
   END dout0[310]
   PIN dout0[311]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1156.68 582.76 1157.06 583.82 ;
      END
   END dout0[311]
   PIN dout0[312]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1158.04 582.76 1158.42 583.82 ;
      END
   END dout0[312]
   PIN dout0[313]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1161.44 582.76 1161.82 583.82 ;
      END
   END dout0[313]
   PIN dout0[314]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1163.48 582.76 1163.86 583.82 ;
      END
   END dout0[314]
   PIN dout0[315]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1167.56 582.76 1167.94 583.82 ;
      END
   END dout0[315]
   PIN dout0[316]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1168.24 582.76 1168.62 583.82 ;
      END
   END dout0[316]
   PIN dout0[317]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1172.32 582.76 1172.7 583.82 ;
      END
   END dout0[317]
   PIN dout0[318]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1173.0 582.76 1173.38 583.82 ;
      END
   END dout0[318]
   PIN dout0[319]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1176.4 582.76 1176.78 583.82 ;
      END
   END dout0[319]
   PIN dout0[320]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1177.76 582.76 1178.14 583.82 ;
      END
   END dout0[320]
   PIN dout0[321]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1182.52 582.76 1182.9 583.82 ;
      END
   END dout0[321]
   PIN dout0[322]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1183.88 582.76 1184.26 583.82 ;
      END
   END dout0[322]
   PIN dout0[323]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1186.6 582.76 1186.98 583.82 ;
      END
   END dout0[323]
   PIN dout0[324]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1187.96 582.76 1188.34 583.82 ;
      END
   END dout0[324]
   PIN dout0[325]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1192.04 582.76 1192.42 583.82 ;
      END
   END dout0[325]
   PIN dout0[326]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1192.72 582.76 1193.1 583.82 ;
      END
   END dout0[326]
   PIN dout0[327]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1197.48 582.76 1197.86 583.82 ;
      END
   END dout0[327]
   PIN dout0[328]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1198.16 582.76 1198.54 583.82 ;
      END
   END dout0[328]
   PIN dout0[329]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1202.24 582.76 1202.62 583.82 ;
      END
   END dout0[329]
   PIN dout0[330]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1203.6 582.76 1203.98 583.82 ;
      END
   END dout0[330]
   PIN dout0[331]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1206.32 582.76 1206.7 583.82 ;
      END
   END dout0[331]
   PIN dout0[332]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1207.68 582.76 1208.06 583.82 ;
      END
   END dout0[332]
   PIN dout0[333]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1211.76 582.76 1212.14 583.82 ;
      END
   END dout0[333]
   PIN dout0[334]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1213.12 582.76 1213.5 583.82 ;
      END
   END dout0[334]
   PIN dout0[335]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1216.52 582.76 1216.9 583.82 ;
      END
   END dout0[335]
   PIN dout0[336]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  1218.56 582.76 1218.94 583.82 ;
      END
   END dout0[336]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.4 3.4 2538.82 5.14 ;
         LAYER met3 ;
         RECT  3.4 578.68 2538.82 580.42 ;
         LAYER met4 ;
         RECT  3.4 3.4 5.14 580.42 ;
         LAYER met4 ;
         RECT  2537.08 3.4 2538.82 580.42 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  2540.48 0.0 2542.22 583.82 ;
         LAYER met3 ;
         RECT  0.0 0.0 2542.22 1.74 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 583.82 ;
         LAYER met3 ;
         RECT  0.0 582.08 2542.22 583.82 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 2541.6 583.2 ;
   LAYER  met2 ;
      RECT  0.62 0.62 2541.6 583.2 ;
   LAYER  met3 ;
      RECT  1.66 279.56 2541.6 281.14 ;
      RECT  0.62 281.82 1.66 287.72 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 279.56 ;
      RECT  2.8 5.74 2539.42 279.56 ;
      RECT  2539.42 2.8 2541.6 5.74 ;
      RECT  2539.42 5.74 2541.6 279.56 ;
      RECT  1.66 281.14 2.8 578.08 ;
      RECT  1.66 578.08 2.8 581.02 ;
      RECT  2.8 281.14 2539.42 578.08 ;
      RECT  2539.42 281.14 2541.6 578.08 ;
      RECT  2539.42 578.08 2541.6 581.02 ;
      RECT  0.62 2.34 1.66 279.56 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 2539.42 2.8 ;
      RECT  2539.42 2.34 2541.6 2.8 ;
      RECT  0.62 289.3 1.66 581.48 ;
      RECT  1.66 581.02 2.8 581.48 ;
      RECT  2.8 581.02 2539.42 581.48 ;
      RECT  2539.42 581.02 2541.6 581.48 ;
   LAYER  met4 ;
      RECT  557.22 0.62 561.76 1.66 ;
      RECT  563.34 0.62 567.88 1.66 ;
      RECT  569.46 0.62 572.64 1.66 ;
      RECT  574.22 0.62 579.44 1.66 ;
      RECT  581.02 0.62 585.56 1.66 ;
      RECT  587.14 0.62 591.0 1.66 ;
      RECT  592.58 0.62 597.12 1.66 ;
      RECT  598.7 0.62 603.24 1.66 ;
      RECT  604.82 0.62 608.68 1.66 ;
      RECT  610.26 0.62 614.12 1.66 ;
      RECT  615.7 0.62 620.24 1.66 ;
      RECT  621.82 0.62 625.68 1.66 ;
      RECT  627.26 0.62 632.48 1.66 ;
      RECT  634.06 0.62 637.92 1.66 ;
      RECT  639.5 0.62 644.04 1.66 ;
      RECT  645.62 0.62 649.48 1.66 ;
      RECT  651.06 0.62 655.6 1.66 ;
      RECT  657.18 0.62 661.04 1.66 ;
      RECT  662.62 0.62 666.48 1.66 ;
      RECT  668.06 0.62 671.92 1.66 ;
      RECT  673.5 0.62 678.04 1.66 ;
      RECT  679.62 0.62 684.16 1.66 ;
      RECT  685.74 0.62 689.6 1.66 ;
      RECT  691.18 0.62 695.72 1.66 ;
      RECT  697.3 0.62 701.16 1.66 ;
      RECT  702.74 0.62 707.28 1.66 ;
      RECT  708.86 0.62 714.08 1.66 ;
      RECT  715.66 0.62 719.52 1.66 ;
      RECT  721.1 0.62 724.96 1.66 ;
      RECT  726.54 0.62 731.76 1.66 ;
      RECT  733.34 0.62 737.2 1.66 ;
      RECT  738.78 0.62 742.64 1.66 ;
      RECT  744.22 0.62 748.08 1.66 ;
      RECT  749.66 0.62 754.2 1.66 ;
      RECT  755.78 0.62 760.32 1.66 ;
      RECT  761.9 0.62 766.44 1.66 ;
      RECT  768.02 0.62 771.2 1.66 ;
      RECT  772.78 0.62 778.0 1.66 ;
      RECT  779.58 0.62 784.12 1.66 ;
      RECT  785.7 0.62 789.56 1.66 ;
      RECT  791.14 0.62 795.68 1.66 ;
      RECT  797.26 0.62 801.12 1.66 ;
      RECT  802.7 0.62 806.56 1.66 ;
      RECT  808.14 0.62 813.36 1.66 ;
      RECT  814.94 0.62 818.12 1.66 ;
      RECT  819.7 0.62 824.92 1.66 ;
      RECT  826.5 0.62 829.68 1.66 ;
      RECT  831.26 0.62 836.48 1.66 ;
      RECT  838.06 0.62 842.6 1.66 ;
      RECT  844.18 0.62 848.04 1.66 ;
      RECT  849.62 0.62 853.48 1.66 ;
      RECT  855.06 0.62 859.6 1.66 ;
      RECT  861.18 0.62 865.72 1.66 ;
      RECT  867.3 0.62 871.84 1.66 ;
      RECT  873.42 0.62 877.28 1.66 ;
      RECT  878.86 0.62 882.72 1.66 ;
      RECT  884.3 0.62 888.84 1.66 ;
      RECT  890.42 0.62 894.28 1.66 ;
      RECT  895.86 0.62 900.4 1.66 ;
      RECT  901.98 0.62 906.52 1.66 ;
      RECT  908.1 0.62 911.96 1.66 ;
      RECT  913.54 0.62 917.4 1.66 ;
      RECT  918.98 0.62 924.2 1.66 ;
      RECT  925.78 0.62 928.96 1.66 ;
      RECT  930.54 0.62 935.08 1.66 ;
      RECT  936.66 0.62 941.2 1.66 ;
      RECT  942.78 0.62 947.32 1.66 ;
      RECT  948.9 0.62 952.76 1.66 ;
      RECT  954.34 0.62 958.88 1.66 ;
      RECT  960.46 0.62 965.0 1.66 ;
      RECT  966.58 0.62 969.76 1.66 ;
      RECT  971.34 0.62 975.88 1.66 ;
      RECT  977.46 0.62 982.68 1.66 ;
      RECT  984.26 0.62 987.44 1.66 ;
      RECT  989.02 0.62 994.24 1.66 ;
      RECT  995.82 0.62 1000.36 1.66 ;
      RECT  1001.94 0.62 1005.8 1.66 ;
      RECT  1007.38 0.62 1011.24 1.66 ;
      RECT  1012.82 0.62 1017.36 1.66 ;
      RECT  1018.94 0.62 1022.8 1.66 ;
      RECT  1024.38 0.62 1029.6 1.66 ;
      RECT  1031.18 0.62 1035.04 1.66 ;
      RECT  1036.62 0.62 1041.16 1.66 ;
      RECT  1042.74 0.62 1046.6 1.66 ;
      RECT  1048.18 0.62 1052.72 1.66 ;
      RECT  1054.3 0.62 1058.16 1.66 ;
      RECT  1059.74 0.62 1064.28 1.66 ;
      RECT  1065.86 0.62 1070.4 1.66 ;
      RECT  1071.98 0.62 1075.84 1.66 ;
      RECT  1077.42 0.62 1081.28 1.66 ;
      RECT  1082.86 0.62 1087.4 1.66 ;
      RECT  1088.98 0.62 1093.52 1.66 ;
      RECT  1095.1 0.62 1098.28 1.66 ;
      RECT  1099.86 0.62 1105.08 1.66 ;
      RECT  1106.66 0.62 1111.2 1.66 ;
      RECT  1112.78 0.62 1115.96 1.66 ;
      RECT  1117.54 0.62 1122.76 1.66 ;
      RECT  1124.34 0.62 1128.2 1.66 ;
      RECT  1129.78 0.62 1133.64 1.66 ;
      RECT  1135.22 0.62 1139.76 1.66 ;
      RECT  1141.34 0.62 1145.88 1.66 ;
      RECT  1147.46 0.62 1152.0 1.66 ;
      RECT  1153.58 0.62 1157.44 1.66 ;
      RECT  1159.02 0.62 1162.88 1.66 ;
      RECT  1164.46 0.62 1169.0 1.66 ;
      RECT  1170.58 0.62 1174.44 1.66 ;
      RECT  1176.02 0.62 1181.24 1.66 ;
      RECT  1182.82 0.62 1186.68 1.66 ;
      RECT  1188.26 0.62 1192.8 1.66 ;
      RECT  1194.38 0.62 1198.24 1.66 ;
      RECT  1199.82 0.62 1204.36 1.66 ;
      RECT  1205.94 0.62 1210.48 1.66 ;
      RECT  1212.06 0.62 1215.92 1.66 ;
      RECT  1217.5 0.62 1222.04 1.66 ;
      RECT  1223.62 0.62 1226.8 1.66 ;
      RECT  1228.38 0.62 1233.6 1.66 ;
      RECT  1235.18 0.62 1239.04 1.66 ;
      RECT  1240.62 0.62 1245.16 1.66 ;
      RECT  1246.74 0.62 1250.6 1.66 ;
      RECT  1252.18 0.62 1256.72 1.66 ;
      RECT  1258.3 0.62 1262.84 1.66 ;
      RECT  1264.42 0.62 1267.6 1.66 ;
      RECT  1269.18 0.62 1274.4 1.66 ;
      RECT  1275.98 0.62 1280.52 1.66 ;
      RECT  1282.1 0.62 1285.96 1.66 ;
      RECT  1287.54 0.62 1291.4 1.66 ;
      RECT  1292.98 0.62 1297.52 1.66 ;
      RECT  1299.1 0.62 1302.96 1.66 ;
      RECT  1304.54 0.62 1309.08 1.66 ;
      RECT  1310.66 0.62 1315.2 1.66 ;
      RECT  1316.78 0.62 1320.64 1.66 ;
      RECT  1322.22 0.62 1327.44 1.66 ;
      RECT  1329.02 0.62 1332.2 1.66 ;
      RECT  1333.78 0.62 1339.0 1.66 ;
      RECT  1340.58 0.62 1344.44 1.66 ;
      RECT  1346.02 0.62 1350.56 1.66 ;
      RECT  1352.14 0.62 1355.32 1.66 ;
      RECT  1356.9 0.62 1362.12 1.66 ;
      RECT  1363.7 0.62 1367.56 1.66 ;
      RECT  1369.14 0.62 1373.0 1.66 ;
      RECT  1374.58 0.62 1379.12 1.66 ;
      RECT  1380.7 0.62 1385.24 1.66 ;
      RECT  1386.82 0.62 1391.36 1.66 ;
      RECT  1392.94 0.62 1397.48 1.66 ;
      RECT  1399.06 0.62 1402.92 1.66 ;
      RECT  1404.5 0.62 1409.04 1.66 ;
      RECT  1410.62 0.62 1414.48 1.66 ;
      RECT  1416.06 0.62 1420.6 1.66 ;
      RECT  1422.18 0.62 1426.72 1.66 ;
      RECT  1428.3 0.62 1431.48 1.66 ;
      RECT  1433.06 0.62 1438.28 1.66 ;
      RECT  1439.86 0.62 1443.72 1.66 ;
      RECT  1445.3 0.62 1449.84 1.66 ;
      RECT  1451.42 0.62 1455.28 1.66 ;
      RECT  1456.86 0.62 1461.4 1.66 ;
      RECT  1462.98 0.62 1467.52 1.66 ;
      RECT  1469.1 0.62 1472.96 1.66 ;
      RECT  1474.54 0.62 1478.4 1.66 ;
      RECT  1479.98 0.62 1483.84 1.66 ;
      RECT  1485.42 0.62 1490.64 1.66 ;
      RECT  1492.22 0.62 1496.08 1.66 ;
      RECT  1497.66 0.62 1502.2 1.66 ;
      RECT  1503.78 0.62 1507.64 1.66 ;
      RECT  1509.22 0.62 1513.76 1.66 ;
      RECT  1515.34 0.62 1519.2 1.66 ;
      RECT  1520.78 0.62 1524.64 1.66 ;
      RECT  1526.22 0.62 1530.76 1.66 ;
      RECT  1532.34 0.62 1536.88 1.66 ;
      RECT  1538.46 0.62 1542.32 1.66 ;
      RECT  1543.9 0.62 1548.44 1.66 ;
      RECT  1550.02 0.62 1553.88 1.66 ;
      RECT  1555.46 0.62 1560.0 1.66 ;
      RECT  1561.58 0.62 1566.12 1.66 ;
      RECT  1567.7 0.62 1572.24 1.66 ;
      RECT  1573.82 0.62 1578.36 1.66 ;
      RECT  1579.94 0.62 1583.12 1.66 ;
      RECT  1584.7 0.62 1589.92 1.66 ;
      RECT  1591.5 0.62 1595.36 1.66 ;
      RECT  1596.94 0.62 1600.8 1.66 ;
      RECT  1602.38 0.62 1607.6 1.66 ;
      RECT  1609.18 0.62 1612.36 1.66 ;
      RECT  1613.94 0.62 1619.16 1.66 ;
      RECT  1620.74 0.62 1625.28 1.66 ;
      RECT  1626.86 0.62 1630.72 1.66 ;
      RECT  1632.3 0.62 1636.16 1.66 ;
      RECT  1637.74 0.62 1642.28 1.66 ;
      RECT  1643.86 0.62 1647.72 1.66 ;
      RECT  1649.3 0.62 1653.84 1.66 ;
      RECT  1655.42 0.62 1659.96 1.66 ;
      RECT  1661.54 0.62 1664.72 1.66 ;
      RECT  1666.3 0.62 1671.52 1.66 ;
      RECT  1673.1 0.62 1676.96 1.66 ;
      RECT  1678.54 0.62 1683.08 1.66 ;
      RECT  1684.66 0.62 1689.2 1.66 ;
      RECT  1690.78 0.62 1694.64 1.66 ;
      RECT  1696.22 0.62 1700.76 1.66 ;
      RECT  1702.34 0.62 1706.2 1.66 ;
      RECT  1707.78 0.62 1712.32 1.66 ;
      RECT  1713.9 0.62 1718.44 1.66 ;
      RECT  1720.02 0.62 1724.56 1.66 ;
      RECT  1726.14 0.62 1730.0 1.66 ;
      RECT  1731.58 0.62 1736.12 1.66 ;
      RECT  1737.7 0.62 1740.88 1.66 ;
      RECT  1742.46 0.62 1747.68 1.66 ;
      RECT  1749.26 0.62 1752.44 1.66 ;
      RECT  1754.02 0.62 1759.24 1.66 ;
      RECT  1760.82 0.62 1764.68 1.66 ;
      RECT  1766.26 0.62 1770.8 1.66 ;
      RECT  1772.38 0.62 1776.24 1.66 ;
      RECT  1777.82 0.62 1782.36 1.66 ;
      RECT  1783.94 0.62 1787.8 1.66 ;
      RECT  1789.38 0.62 1794.6 1.66 ;
      RECT  1796.18 0.62 1799.36 1.66 ;
      RECT  1800.94 0.62 1805.48 1.66 ;
      RECT  1807.06 0.62 1811.6 1.66 ;
      RECT  1813.18 0.62 1817.04 1.66 ;
      RECT  1818.62 0.62 1822.48 1.66 ;
      RECT  1824.06 0.62 1829.28 1.66 ;
      RECT  1830.86 0.62 1835.4 1.66 ;
      RECT  1836.98 0.62 1840.84 1.66 ;
      RECT  1842.42 0.62 1846.28 1.66 ;
      RECT  1847.86 0.62 1852.4 1.66 ;
      RECT  1853.98 0.62 1858.52 1.66 ;
      RECT  1860.1 0.62 1863.28 1.66 ;
      RECT  1864.86 0.62 1870.08 1.66 ;
      RECT  1871.66 0.62 1876.2 1.66 ;
      RECT  1877.78 0.62 1880.96 1.66 ;
      RECT  1882.54 0.62 1887.76 1.66 ;
      RECT  1889.34 0.62 1892.52 1.66 ;
      RECT  1894.1 0.62 1899.32 1.66 ;
      RECT  1900.9 0.62 1905.44 1.66 ;
      RECT  1907.02 0.62 1910.88 1.66 ;
      RECT  1912.46 0.62 1916.32 1.66 ;
      RECT  1917.9 0.62 1921.76 1.66 ;
      RECT  1923.34 0.62 1927.88 1.66 ;
      RECT  1929.46 0.62 1934.0 1.66 ;
      RECT  1935.58 0.62 1939.44 1.66 ;
      RECT  1941.02 0.62 1945.56 1.66 ;
      RECT  1947.14 0.62 1951.0 1.66 ;
      RECT  1952.58 0.62 1957.12 1.66 ;
      RECT  1958.7 0.62 1962.56 1.66 ;
      RECT  1964.14 0.62 1968.68 1.66 ;
      RECT  1970.26 0.62 1975.48 1.66 ;
      RECT  1977.06 0.62 1980.24 1.66 ;
      RECT  1981.82 0.62 1986.36 1.66 ;
      RECT  1987.94 0.62 1992.48 1.66 ;
      RECT  1994.06 0.62 1997.92 1.66 ;
      RECT  1999.5 0.62 2004.04 1.66 ;
      RECT  2005.62 0.62 2010.16 1.66 ;
      RECT  2011.74 0.62 2016.28 1.66 ;
      RECT  2017.86 0.62 2022.4 1.66 ;
      RECT  2023.98 0.62 2027.84 1.66 ;
      RECT  2029.42 0.62 2033.96 1.66 ;
      RECT  2035.54 0.62 2039.4 1.66 ;
      RECT  2040.98 0.62 2045.52 1.66 ;
      RECT  2047.1 0.62 2050.28 1.66 ;
      RECT  2051.86 0.62 2057.08 1.66 ;
      RECT  2058.66 0.62 2061.84 1.66 ;
      RECT  2063.42 0.62 2068.64 1.66 ;
      RECT  2070.22 0.62 2074.08 1.66 ;
      RECT  2075.66 0.62 2080.2 1.66 ;
      RECT  2081.78 0.62 2085.64 1.66 ;
      RECT  2087.22 0.62 2091.76 1.66 ;
      RECT  2093.34 0.62 2097.2 1.66 ;
      RECT  2098.78 0.62 2103.32 1.66 ;
      RECT  2104.9 0.62 2108.76 1.66 ;
      RECT  2110.34 0.62 2115.56 1.66 ;
      RECT  2117.14 0.62 2121.68 1.66 ;
      RECT  2123.26 0.62 2127.12 1.66 ;
      RECT  2128.7 0.62 2132.56 1.66 ;
      RECT  2134.14 0.62 2138.68 1.66 ;
      RECT  2140.26 0.62 2144.12 1.66 ;
      RECT  2145.7 0.62 2150.24 1.66 ;
      RECT  2151.82 0.62 2155.68 1.66 ;
      RECT  2157.26 0.62 2161.8 1.66 ;
      RECT  2163.38 0.62 2167.24 1.66 ;
      RECT  2168.82 0.62 2173.36 1.66 ;
      RECT  2174.94 0.62 2179.48 1.66 ;
      RECT  2181.06 0.62 2184.92 1.66 ;
      RECT  2186.5 0.62 2191.04 1.66 ;
      RECT  2192.62 0.62 2196.48 1.66 ;
      RECT  2198.06 0.62 2203.28 1.66 ;
      RECT  2204.86 0.62 2208.04 1.66 ;
      RECT  2209.62 0.62 2214.16 1.66 ;
      RECT  2215.74 0.62 2219.6 1.66 ;
      RECT  2221.18 0.62 2225.72 1.66 ;
      RECT  2227.3 0.62 2232.52 1.66 ;
      RECT  2234.1 0.62 2237.28 1.66 ;
      RECT  2238.86 0.62 2244.08 1.66 ;
      RECT  2245.66 0.62 2248.84 1.66 ;
      RECT  2250.42 0.62 2255.64 1.66 ;
      RECT  2257.22 0.62 2260.4 1.66 ;
      RECT  2261.98 0.62 2267.2 1.66 ;
      RECT  2268.78 0.62 2272.64 1.66 ;
      RECT  2274.22 0.62 2278.76 1.66 ;
      RECT  2280.34 0.62 2284.88 1.66 ;
      RECT  2286.46 0.62 2290.32 1.66 ;
      RECT  2291.9 0.62 2296.44 1.66 ;
      RECT  2298.02 0.62 2302.56 1.66 ;
      RECT  2304.14 0.62 2308.0 1.66 ;
      RECT  2309.58 0.62 2314.12 1.66 ;
      RECT  2315.7 0.62 2319.56 1.66 ;
      RECT  2321.14 0.62 2325.68 1.66 ;
      RECT  2327.26 0.62 2331.12 1.66 ;
      RECT  2332.7 0.62 2337.24 1.66 ;
      RECT  2338.82 0.62 2343.36 1.66 ;
      RECT  2344.94 0.62 2348.12 1.66 ;
      RECT  2349.7 0.62 2354.92 1.66 ;
      RECT  2356.5 0.62 2359.68 1.66 ;
      RECT  2361.26 0.62 2365.8 1.66 ;
      RECT  2367.38 0.62 2371.92 1.66 ;
      RECT  2373.5 0.62 2377.36 1.66 ;
      RECT  2378.94 0.62 2384.16 1.66 ;
      RECT  2385.74 0.62 2390.28 1.66 ;
      RECT  2391.86 0.62 2395.72 1.66 ;
      RECT  2397.3 0.62 2401.16 1.66 ;
      RECT  2402.74 0.62 2407.28 1.66 ;
      RECT  2408.86 0.62 2412.72 1.66 ;
      RECT  2414.3 0.62 2418.16 1.66 ;
      RECT  2419.74 0.62 2424.28 1.66 ;
      RECT  2425.86 0.62 2430.4 1.66 ;
      RECT  2431.98 0.62 2436.52 1.66 ;
      RECT  2438.1 0.62 2441.96 1.66 ;
      RECT  2443.54 0.62 2447.4 1.66 ;
      RECT  2448.98 0.62 2454.2 1.66 ;
      RECT  2455.78 0.62 2460.32 1.66 ;
      RECT  2461.9 0.62 2465.76 1.66 ;
      RECT  2467.34 0.62 2471.2 1.66 ;
      RECT  2472.78 0.62 2477.32 1.66 ;
      RECT  2478.9 0.62 2482.76 1.66 ;
      RECT  2484.34 0.62 2488.88 1.66 ;
      RECT  2490.46 0.62 2494.32 1.66 ;
      RECT  2495.9 0.62 2501.12 1.66 ;
      RECT  2502.7 0.62 2505.88 1.66 ;
      RECT  2507.46 0.62 2512.68 1.66 ;
      RECT  2514.26 0.62 2518.8 1.66 ;
      RECT  295.88 1.66 297.46 582.16 ;
      RECT  297.46 1.66 555.64 582.16 ;
      RECT  298.82 582.16 299.28 583.2 ;
      RECT  312.42 0.62 316.28 1.66 ;
      RECT  317.86 0.62 322.4 1.66 ;
      RECT  323.98 0.62 327.84 1.66 ;
      RECT  329.42 0.62 333.96 1.66 ;
      RECT  335.54 0.62 339.4 1.66 ;
      RECT  340.98 0.62 346.2 1.66 ;
      RECT  347.78 0.62 350.96 1.66 ;
      RECT  352.54 0.62 357.76 1.66 ;
      RECT  359.34 0.62 362.52 1.66 ;
      RECT  364.1 0.62 369.32 1.66 ;
      RECT  370.9 0.62 375.44 1.66 ;
      RECT  377.02 0.62 380.88 1.66 ;
      RECT  382.46 0.62 386.32 1.66 ;
      RECT  387.9 0.62 392.44 1.66 ;
      RECT  394.02 0.62 397.88 1.66 ;
      RECT  399.46 0.62 404.68 1.66 ;
      RECT  406.26 0.62 409.44 1.66 ;
      RECT  411.02 0.62 416.24 1.66 ;
      RECT  417.82 0.62 421.0 1.66 ;
      RECT  422.58 0.62 427.8 1.66 ;
      RECT  429.38 0.62 432.56 1.66 ;
      RECT  434.14 0.62 439.36 1.66 ;
      RECT  440.94 0.62 444.8 1.66 ;
      RECT  446.38 0.62 450.92 1.66 ;
      RECT  452.5 0.62 456.36 1.66 ;
      RECT  457.94 0.62 462.48 1.66 ;
      RECT  464.06 0.62 468.6 1.66 ;
      RECT  470.18 0.62 474.72 1.66 ;
      RECT  476.3 0.62 480.16 1.66 ;
      RECT  481.74 0.62 486.28 1.66 ;
      RECT  487.86 0.62 491.04 1.66 ;
      RECT  492.62 0.62 497.84 1.66 ;
      RECT  499.42 0.62 502.6 1.66 ;
      RECT  504.18 0.62 509.4 1.66 ;
      RECT  510.98 0.62 514.84 1.66 ;
      RECT  516.42 0.62 520.28 1.66 ;
      RECT  521.86 0.62 527.08 1.66 ;
      RECT  528.66 0.62 533.2 1.66 ;
      RECT  534.78 0.62 538.64 1.66 ;
      RECT  540.22 0.62 544.08 1.66 ;
      RECT  545.66 0.62 549.52 1.66 ;
      RECT  551.1 0.62 555.64 1.66 ;
      RECT  2520.38 0.62 2524.24 1.66 ;
      RECT  303.58 582.16 377.48 583.2 ;
      RECT  379.06 582.16 381.56 583.2 ;
      RECT  384.5 582.16 385.64 583.2 ;
      RECT  387.22 582.16 387.68 583.2 ;
      RECT  389.26 582.16 391.08 583.2 ;
      RECT  392.66 582.16 393.12 583.2 ;
      RECT  394.7 582.16 395.84 583.2 ;
      RECT  398.78 582.16 401.96 583.2 ;
      RECT  404.22 582.16 406.72 583.2 ;
      RECT  408.98 582.16 410.8 583.2 ;
      RECT  413.74 582.16 416.92 583.2 ;
      RECT  419.86 582.16 421.68 583.2 ;
      RECT  423.94 582.16 425.76 583.2 ;
      RECT  428.7 582.16 431.88 583.2 ;
      RECT  434.82 582.16 435.96 583.2 ;
      RECT  438.9 582.16 441.4 583.2 ;
      RECT  444.34 582.16 446.84 583.2 ;
      RECT  449.1 582.16 450.92 583.2 ;
      RECT  453.86 582.16 455.68 583.2 ;
      RECT  458.62 582.16 461.8 583.2 ;
      RECT  464.06 582.16 466.56 583.2 ;
      RECT  468.82 582.16 470.64 583.2 ;
      RECT  473.58 582.16 476.76 583.2 ;
      RECT  479.7 582.16 481.52 583.2 ;
      RECT  484.46 582.16 486.96 583.2 ;
      RECT  489.22 582.16 491.04 583.2 ;
      RECT  492.62 582.16 493.08 583.2 ;
      RECT  494.66 582.16 495.8 583.2 ;
      RECT  498.74 582.16 501.24 583.2 ;
      RECT  504.18 582.16 506.68 583.2 ;
      RECT  508.94 582.16 510.76 583.2 ;
      RECT  512.34 582.16 512.8 583.2 ;
      RECT  514.38 582.16 516.88 583.2 ;
      RECT  519.82 582.16 520.96 583.2 ;
      RECT  523.9 582.16 525.72 583.2 ;
      RECT  528.66 582.16 531.16 583.2 ;
      RECT  534.1 582.16 535.92 583.2 ;
      RECT  537.5 582.16 537.96 583.2 ;
      RECT  539.54 582.16 540.68 583.2 ;
      RECT  543.62 582.16 546.8 583.2 ;
      RECT  549.06 582.16 550.88 583.2 ;
      RECT  553.82 582.16 555.64 583.2 ;
      RECT  555.64 1.66 557.22 582.16 ;
      RECT  557.22 1.66 558.58 582.16 ;
      RECT  558.58 582.16 561.08 583.2 ;
      RECT  564.02 582.16 565.84 583.2 ;
      RECT  568.78 582.16 571.96 583.2 ;
      RECT  574.22 582.16 576.72 583.2 ;
      RECT  579.66 582.16 580.8 583.2 ;
      RECT  583.74 582.16 586.92 583.2 ;
      RECT  589.18 582.16 591.0 583.2 ;
      RECT  593.94 582.16 595.76 583.2 ;
      RECT  597.34 582.16 597.8 583.2 ;
      RECT  599.38 582.16 601.88 583.2 ;
      RECT  604.14 582.16 606.64 583.2 ;
      RECT  608.9 582.16 610.72 583.2 ;
      RECT  613.66 582.16 616.84 583.2 ;
      RECT  619.78 582.16 621.6 583.2 ;
      RECT  624.54 582.16 626.36 583.2 ;
      RECT  628.62 582.16 631.12 583.2 ;
      RECT  634.06 582.16 635.88 583.2 ;
      RECT  637.46 582.16 637.92 583.2 ;
      RECT  639.5 582.16 640.64 583.2 ;
      RECT  642.22 582.16 642.68 583.2 ;
      RECT  644.26 582.16 646.08 583.2 ;
      RECT  649.02 582.16 650.84 583.2 ;
      RECT  653.78 582.16 656.96 583.2 ;
      RECT  659.22 582.16 661.72 583.2 ;
      RECT  664.66 582.16 666.48 583.2 ;
      RECT  668.74 582.16 671.92 583.2 ;
      RECT  674.86 582.16 676.68 583.2 ;
      RECT  679.62 582.16 680.76 583.2 ;
      RECT  683.7 582.16 686.2 583.2 ;
      RECT  689.14 582.16 690.96 583.2 ;
      RECT  693.9 582.16 696.4 583.2 ;
      RECT  699.34 582.16 701.84 583.2 ;
      RECT  704.1 582.16 705.92 583.2 ;
      RECT  708.86 582.16 710.68 583.2 ;
      RECT  713.62 582.16 716.8 583.2 ;
      RECT  719.06 582.16 720.88 583.2 ;
      RECT  723.82 582.16 725.64 583.2 ;
      RECT  727.22 582.16 727.68 583.2 ;
      RECT  729.26 582.16 731.76 583.2 ;
      RECT  734.02 582.16 735.84 583.2 ;
      RECT  738.78 582.16 741.96 583.2 ;
      RECT  744.22 582.16 746.04 583.2 ;
      RECT  748.98 582.16 751.48 583.2 ;
      RECT  753.74 582.16 756.24 583.2 ;
      RECT  757.82 582.16 758.28 583.2 ;
      RECT  759.86 582.16 761.68 583.2 ;
      RECT  763.94 582.16 765.76 583.2 ;
      RECT  768.7 582.16 771.2 583.2 ;
      RECT  774.14 582.16 775.96 583.2 ;
      RECT  778.9 582.16 781.4 583.2 ;
      RECT  783.66 582.16 786.16 583.2 ;
      RECT  789.1 582.16 790.92 583.2 ;
      RECT  793.86 582.16 795.68 583.2 ;
      RECT  798.62 582.16 801.8 583.2 ;
      RECT  804.06 582.16 805.88 583.2 ;
      RECT  808.82 582.16 810.64 583.2 ;
      RECT  812.22 582.16 812.68 583.2 ;
      RECT  814.26 582.16 816.08 583.2 ;
      RECT  817.66 582.16 818.12 583.2 ;
      RECT  819.7 582.16 821.52 583.2 ;
      RECT  823.78 582.16 826.96 583.2 ;
      RECT  829.22 582.16 831.04 583.2 ;
      RECT  833.98 582.16 835.8 583.2 ;
      RECT  838.74 582.16 841.92 583.2 ;
      RECT  844.18 582.16 846.0 583.2 ;
      RECT  848.94 582.16 850.76 583.2 ;
      RECT  853.7 582.16 856.88 583.2 ;
      RECT  859.82 582.16 861.64 583.2 ;
      RECT  863.9 582.16 865.72 583.2 ;
      RECT  868.66 582.16 871.16 583.2 ;
      RECT  874.1 582.16 876.6 583.2 ;
      RECT  878.86 582.16 880.68 583.2 ;
      RECT  882.26 582.16 882.72 583.2 ;
      RECT  884.3 582.16 886.8 583.2 ;
      RECT  889.06 582.16 890.88 583.2 ;
      RECT  893.82 582.16 895.64 583.2 ;
      RECT  897.22 582.16 897.68 583.2 ;
      RECT  899.26 582.16 901.08 583.2 ;
      RECT  904.02 582.16 905.84 583.2 ;
      RECT  908.78 582.16 911.28 583.2 ;
      RECT  914.22 582.16 916.04 583.2 ;
      RECT  918.98 582.16 920.8 583.2 ;
      RECT  922.38 582.16 922.84 583.2 ;
      RECT  924.42 582.16 926.92 583.2 ;
      RECT  929.18 582.16 931.0 583.2 ;
      RECT  933.94 582.16 935.76 583.2 ;
      RECT  938.7 582.16 941.2 583.2 ;
      RECT  944.14 582.16 946.64 583.2 ;
      RECT  948.9 582.16 951.4 583.2 ;
      RECT  953.66 582.16 956.84 583.2 ;
      RECT  959.78 582.16 960.92 583.2 ;
      RECT  962.5 582.16 962.96 583.2 ;
      RECT  964.54 582.16 966.36 583.2 ;
      RECT  969.3 582.16 971.12 583.2 ;
      RECT  974.06 582.16 975.88 583.2 ;
      RECT  978.82 582.16 981.32 583.2 ;
      RECT  984.26 582.16 986.08 583.2 ;
      RECT  989.02 582.16 990.84 583.2 ;
      RECT  993.78 582.16 996.96 583.2 ;
      RECT  999.22 582.16 1001.04 583.2 ;
      RECT  1003.98 582.16 1006.48 583.2 ;
      RECT  1009.42 582.16 1011.92 583.2 ;
      RECT  1014.86 582.16 1016.0 583.2 ;
      RECT  1018.94 582.16 1020.76 583.2 ;
      RECT  1023.7 582.16 1026.88 583.2 ;
      RECT  1029.14 582.16 1031.64 583.2 ;
      RECT  1033.9 582.16 1036.4 583.2 ;
      RECT  1039.34 582.16 1041.16 583.2 ;
      RECT  1042.74 582.16 1043.2 583.2 ;
      RECT  1044.78 582.16 1046.6 583.2 ;
      RECT  1048.86 582.16 1050.68 583.2 ;
      RECT  1052.26 582.16 1052.72 583.2 ;
      RECT  1054.3 582.16 1056.8 583.2 ;
      RECT  1059.06 582.16 1060.88 583.2 ;
      RECT  1063.82 582.16 1066.32 583.2 ;
      RECT  1069.26 582.16 1071.08 583.2 ;
      RECT  1074.02 582.16 1075.84 583.2 ;
      RECT  1077.42 582.16 1077.88 583.2 ;
      RECT  1079.46 582.16 1081.96 583.2 ;
      RECT  1084.9 582.16 1086.72 583.2 ;
      RECT  1088.98 582.16 1090.8 583.2 ;
      RECT  1093.74 582.16 1096.92 583.2 ;
      RECT  1099.18 582.16 1101.68 583.2 ;
      RECT  1104.62 582.16 1106.44 583.2 ;
      RECT  1109.38 582.16 1111.88 583.2 ;
      RECT  1114.14 582.16 1115.96 583.2 ;
      RECT  1117.54 582.16 1118.0 583.2 ;
      RECT  1119.58 582.16 1120.72 583.2 ;
      RECT  1123.66 582.16 1126.16 583.2 ;
      RECT  1129.1 582.16 1130.92 583.2 ;
      RECT  1133.86 582.16 1135.68 583.2 ;
      RECT  1137.26 582.16 1137.72 583.2 ;
      RECT  1139.3 582.16 1141.8 583.2 ;
      RECT  1144.74 582.16 1145.88 583.2 ;
      RECT  1148.82 582.16 1150.64 583.2 ;
      RECT  1153.58 582.16 1156.08 583.2 ;
      RECT  1159.02 582.16 1160.84 583.2 ;
      RECT  1162.42 582.16 1162.88 583.2 ;
      RECT  1164.46 582.16 1166.96 583.2 ;
      RECT  1169.22 582.16 1171.72 583.2 ;
      RECT  1173.98 582.16 1175.8 583.2 ;
      RECT  1178.74 582.16 1181.92 583.2 ;
      RECT  1184.86 582.16 1186.0 583.2 ;
      RECT  1188.94 582.16 1191.44 583.2 ;
      RECT  1193.7 582.16 1196.88 583.2 ;
      RECT  1199.14 582.16 1201.64 583.2 ;
      RECT  1204.58 582.16 1205.72 583.2 ;
      RECT  1208.66 582.16 1211.16 583.2 ;
      RECT  1214.1 582.16 1215.92 583.2 ;
      RECT  1217.5 582.16 1217.96 583.2 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 581.02 5.74 582.16 ;
      RECT  5.74 1.66 295.88 2.8 ;
      RECT  5.74 2.8 295.88 581.02 ;
      RECT  5.74 581.02 295.88 582.16 ;
      RECT  558.58 1.66 2536.48 2.8 ;
      RECT  558.58 2.8 2536.48 581.02 ;
      RECT  558.58 581.02 2536.48 582.16 ;
      RECT  2536.48 1.66 2539.42 2.8 ;
      RECT  2536.48 581.02 2539.42 582.16 ;
      RECT  2525.82 0.62 2539.88 1.66 ;
      RECT  1219.54 582.16 2539.88 583.2 ;
      RECT  2539.42 1.66 2539.88 2.8 ;
      RECT  2539.42 2.8 2539.88 581.02 ;
      RECT  2539.42 581.02 2539.88 582.16 ;
      RECT  2.34 582.16 295.88 583.2 ;
      RECT  2.34 0.62 310.84 1.66 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 581.02 ;
      RECT  2.34 581.02 2.8 582.16 ;
   END
END    sram_336x128
END    LIBRARY
