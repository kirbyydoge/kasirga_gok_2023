`define CTR_BIT     5

`define CNTP_STEP   4
`define CNTZ_STEP   4
`define HMDST_STEP  4