`define MATCH_SLLI_RV32         32'h1013
`define MASK_SLLI_RV32          32'hfe00707f
`define MATCH_SRLI_RV32         32'h5013
`define MASK_SRLI_RV32          32'hfe00707f
`define MATCH_SRAI_RV32         32'h40005013
`define MASK_SRAI_RV32          32'hfe00707f
`define MATCH_FRFLAGS           32'h102073
`define MASK_FRFLAGS            32'hfffff07f
`define MATCH_FSFLAGS           32'h101073
`define MASK_FSFLAGS            32'hfff0707f
`define MATCH_FSFLAGSI          32'h105073
`define MASK_FSFLAGSI           32'hfff0707f
`define MATCH_FRRM              32'h202073
`define MASK_FRRM               32'hfffff07f
`define MATCH_FSRM              32'h201073
`define MASK_FSRM               32'hfff0707f
`define MATCH_FSRMI             32'h205073
`define MASK_FSRMI              32'hfff0707f
`define MATCH_FSCSR             32'h301073
`define MASK_FSCSR              32'hfff0707f
`define MATCH_FRCSR             32'h302073
`define MASK_FRCSR              32'hfffff07f
`define MATCH_RDCYCLE           32'hc0002073
`define MASK_RDCYCLE            32'hfffff07f
`define MATCH_RDTIME            32'hc0102073
`define MASK_RDTIME             32'hfffff07f
`define MATCH_RDINSTRET         32'hc0202073
`define MASK_RDINSTRET          32'hfffff07f
`define MATCH_RDCYCLEH          32'hc8002073
`define MASK_RDCYCLEH           32'hfffff07f
`define MATCH_RDTIMEH           32'hc8102073
`define MASK_RDTIMEH            32'hfffff07f
`define MATCH_RDINSTRETH        32'hc8202073
`define MASK_RDINSTRETH         32'hfffff07f
`define MATCH_SCALL             32'h73
`define MASK_SCALL              32'hffffffff
`define MATCH_SBREAK            32'h100073
`define MASK_SBREAK             32'hffffffff
`define MATCH_BEQ               32'h63
`define MASK_BEQ                32'h707f
`define MATCH_BNE               32'h1063
`define MASK_BNE                32'h707f
`define MATCH_BLT               32'h4063
`define MASK_BLT                32'h707f
`define MATCH_BGE               32'h5063
`define MASK_BGE                32'h707f
`define MATCH_BLTU              32'h6063
`define MASK_BLTU               32'h707f
`define MATCH_BGEU              32'h7063
`define MASK_BGEU               32'h707f
`define MATCH_JALR              32'h67
`define MASK_JALR               32'h707f
`define MATCH_JAL               32'h6f
`define MASK_JAL                32'h7f
`define MATCH_LUI               32'h37
`define MASK_LUI                32'h7f
`define MATCH_AUIPC             32'h17
`define MASK_AUIPC              32'h7f
`define MATCH_ADDI              32'h13
`define MASK_ADDI               32'h707f
`define MATCH_SLLI              32'h1013
`define MASK_SLLI               32'hfc00707f
`define MATCH_SLTI              32'h2013
`define MASK_SLTI               32'h707f
`define MATCH_SLTIU             32'h3013
`define MASK_SLTIU              32'h707f
`define MATCH_XORI              32'h4013
`define MASK_XORI               32'h707f
`define MATCH_SRLI              32'h5013
`define MASK_SRLI               32'hfc00707f
`define MATCH_SRAI              32'h40005013
`define MASK_SRAI               32'hfc00707f
`define MATCH_ORI               32'h6013
`define MASK_ORI                32'h707f
`define MATCH_ANDI              32'h7013
`define MASK_ANDI               32'h707f
`define MATCH_ADD               32'h33
`define MASK_ADD                32'hfe00707f
`define MATCH_SUB               32'h40000033
`define MASK_SUB                32'hfe00707f
`define MATCH_SLL               32'h1033
`define MASK_SLL                32'hfe00707f
`define MATCH_SLT               32'h2033
`define MASK_SLT                32'hfe00707f
`define MATCH_SLTU              32'h3033
`define MASK_SLTU               32'hfe00707f
`define MATCH_XOR               32'h4033
`define MASK_XOR                32'hfe00707f
`define MATCH_SRL               32'h5033
`define MASK_SRL                32'hfe00707f
`define MATCH_SRA               32'h40005033
`define MASK_SRA                32'hfe00707f
`define MATCH_OR                32'h6033
`define MASK_OR                 32'hfe00707f
`define MATCH_AND               32'h7033
`define MASK_AND                32'hfe00707f
`define MATCH_ADDIW             32'h1b
`define MASK_ADDIW              32'h707f
`define MATCH_SLLIW             32'h101b
`define MASK_SLLIW              32'hfe00707f
`define MATCH_SRLIW             32'h501b
`define MASK_SRLIW              32'hfe00707f
`define MATCH_SRAIW             32'h4000501b
`define MASK_SRAIW              32'hfe00707f
`define MATCH_ADDW              32'h3b
`define MASK_ADDW               32'hfe00707f
`define MATCH_SUBW              32'h4000003b
`define MASK_SUBW               32'hfe00707f
`define MATCH_SLLW              32'h103b
`define MASK_SLLW               32'hfe00707f
`define MATCH_SRLW              32'h503b
`define MASK_SRLW               32'hfe00707f
`define MATCH_SRAW              32'h4000503b
`define MASK_SRAW               32'hfe00707f
`define MATCH_LB                32'h3
`define MASK_LB                 32'h707f
`define MATCH_LH                32'h1003
`define MASK_LH                 32'h707f
`define MATCH_LW                32'h2003
`define MASK_LW                 32'h707f
`define MATCH_LD                32'h3003
`define MASK_LD                 32'h707f
`define MATCH_LBU               32'h4003
`define MASK_LBU                32'h707f
`define MATCH_LHU               32'h5003
`define MASK_LHU                32'h707f
`define MATCH_LWU               32'h6003
`define MASK_LWU                32'h707f
`define MATCH_SB                32'h23
`define MASK_SB                 32'h707f
`define MATCH_SH                32'h1023
`define MASK_SH                 32'h707f
`define MATCH_SW                32'h2023
`define MASK_SW                 32'h707f
`define MATCH_SD                32'h3023
`define MASK_SD                 32'h707f
`define MATCH_PAUSE             32'h0100000f
`define MASK_PAUSE              32'hffffffff
`define MATCH_FENCE             32'hf
`define MASK_FENCE              32'h707f
`define MATCH_FENCE_I           32'h100f
`define MASK_FENCE_I            32'h707f
`define MATCH_FENCE_TSO         32'h8330000f
`define MASK_FENCE_TSO          32'hfff0707f
`define MATCH_MUL               32'h2000033
`define MASK_MUL                32'hfe00707f
`define MATCH_MULH              32'h2001033
`define MASK_MULH               32'hfe00707f
`define MATCH_MULHSU            32'h2002033
`define MASK_MULHSU             32'hfe00707f
`define MATCH_MULHU             32'h2003033
`define MASK_MULHU              32'hfe00707f
`define MATCH_DIV               32'h2004033
`define MASK_DIV                32'hfe00707f
`define MATCH_DIVU              32'h2005033
`define MASK_DIVU               32'hfe00707f
`define MATCH_REM               32'h2006033
`define MASK_REM                32'hfe00707f
`define MATCH_REMU              32'h2007033
`define MASK_REMU               32'hfe00707f
`define MATCH_MULW              32'h200003b
`define MASK_MULW               32'hfe00707f
`define MATCH_DIVW              32'h200403b
`define MASK_DIVW               32'hfe00707f
`define MATCH_DIVUW             32'h200503b
`define MASK_DIVUW              32'hfe00707f
`define MATCH_REMW              32'h200603b
`define MASK_REMW               32'hfe00707f
`define MATCH_REMUW             32'h200703b
`define MASK_REMUW              32'hfe00707f
`define MATCH_AMOADD_W          32'h202f
`define MASK_AMOADD_W           32'hf800707f
`define MATCH_AMOXOR_W          32'h2000202f
`define MASK_AMOXOR_W           32'hf800707f
`define MATCH_AMOOR_W           32'h4000202f
`define MASK_AMOOR_W            32'hf800707f
`define MATCH_AMOAND_W          32'h6000202f
`define MASK_AMOAND_W           32'hf800707f
`define MATCH_AMOMIN_W          32'h8000202f
`define MASK_AMOMIN_W           32'hf800707f
`define MATCH_AMOMAX_W          32'ha000202f
`define MASK_AMOMAX_W           32'hf800707f
`define MATCH_AMOMINU_W         32'hc000202f
`define MASK_AMOMINU_W          32'hf800707f
`define MATCH_AMOMAXU_W         32'he000202f
`define MASK_AMOMAXU_W          32'hf800707f
`define MATCH_AMOSWAP_W         32'h800202f
`define MASK_AMOSWAP_W          32'hf800707f
`define MATCH_LR_W              32'h1000202f
`define MASK_LR_W               32'hf9f0707f
`define MATCH_SC_W              32'h1800202f
`define MASK_SC_W               32'hf800707f
`define MATCH_AMOADD_D          32'h302f
`define MASK_AMOADD_D           32'hf800707f
`define MATCH_AMOXOR_D          32'h2000302f
`define MASK_AMOXOR_D           32'hf800707f
`define MATCH_AMOOR_D           32'h4000302f
`define MASK_AMOOR_D            32'hf800707f
`define MATCH_AMOAND_D          32'h6000302f
`define MASK_AMOAND_D           32'hf800707f
`define MATCH_AMOMIN_D          32'h8000302f
`define MASK_AMOMIN_D           32'hf800707f
`define MATCH_AMOMAX_D          32'ha000302f
`define MASK_AMOMAX_D           32'hf800707f
`define MATCH_AMOMINU_D         32'hc000302f
`define MASK_AMOMINU_D          32'hf800707f
`define MATCH_AMOMAXU_D         32'he000302f
`define MASK_AMOMAXU_D          32'hf800707f
`define MATCH_AMOSWAP_D         32'h800302f
`define MASK_AMOSWAP_D          32'hf800707f
`define MATCH_LR_D              32'h1000302f
`define MASK_LR_D               32'hf9f0707f
`define MATCH_SC_D              32'h1800302f
`define MASK_SC_D               32'hf800707f
`define MATCH_ECALL             32'h73
`define MASK_ECALL              32'hffffffff
`define MATCH_EBREAK            32'h100073
`define MASK_EBREAK             32'hffffffff
`define MATCH_URET              32'h200073
`define MASK_URET               32'hffffffff
`define MATCH_SRET              32'h10200073
`define MASK_SRET               32'hffffffff
`define MATCH_HRET              32'h20200073
`define MASK_HRET               32'hffffffff
`define MATCH_MRET              32'h30200073
`define MASK_MRET               32'hffffffff
`define MATCH_DRET              32'h7b200073
`define MASK_DRET               32'hffffffff
`define MATCH_SFENCE_VM         32'h10400073
`define MASK_SFENCE_VM          32'hfff07fff
`define MATCH_SFENCE_VMA        32'h12000073
`define MASK_SFENCE_VMA         32'hfe007fff
`define MATCH_WFI               32'h10500073
`define MASK_WFI                32'hffffffff
`define MATCH_CSRRW             32'h1073
`define MASK_CSRRW              32'h707f
`define MATCH_CSRRS             32'h2073
`define MASK_CSRRS              32'h707f
`define MATCH_CSRRC             32'h3073
`define MASK_CSRRC              32'h707f
`define MATCH_CSRRWI            32'h5073
`define MASK_CSRRWI             32'h707f
`define MATCH_CSRRSI            32'h6073
`define MASK_CSRRSI             32'h707f
`define MATCH_CSRRCI            32'h7073
`define MASK_CSRRCI             32'h707f
`define MATCH_FADD_S            32'h53
`define MASK_FADD_S             32'hfe00007f
`define MATCH_FSUB_S            32'h8000053
`define MASK_FSUB_S             32'hfe00007f
`define MATCH_FMUL_S            32'h10000053
`define MASK_FMUL_S             32'hfe00007f
`define MATCH_FDIV_S            32'h18000053
`define MASK_FDIV_S             32'hfe00007f
`define MATCH_FSGNJ_S           32'h20000053
`define MASK_FSGNJ_S            32'hfe00707f
`define MATCH_FSGNJN_S          32'h20001053
`define MASK_FSGNJN_S           32'hfe00707f
`define MATCH_FSGNJX_S          32'h20002053
`define MASK_FSGNJX_S           32'hfe00707f
`define MATCH_FMIN_S            32'h28000053
`define MASK_FMIN_S             32'hfe00707f
`define MATCH_FMAX_S            32'h28001053
`define MASK_FMAX_S             32'hfe00707f
`define MATCH_FSQRT_S           32'h58000053
`define MASK_FSQRT_S            32'hfff0007f
`define MATCH_FADD_D            32'h2000053
`define MASK_FADD_D             32'hfe00007f
`define MATCH_FSUB_D            32'ha000053
`define MASK_FSUB_D             32'hfe00007f
`define MATCH_FMUL_D            32'h12000053
`define MASK_FMUL_D             32'hfe00007f
`define MATCH_FDIV_D            32'h1a000053
`define MASK_FDIV_D             32'hfe00007f
`define MATCH_FSGNJ_D           32'h22000053
`define MASK_FSGNJ_D            32'hfe00707f
`define MATCH_FSGNJN_D          32'h22001053
`define MASK_FSGNJN_D           32'hfe00707f
`define MATCH_FSGNJX_D          32'h22002053
`define MASK_FSGNJX_D           32'hfe00707f
`define MATCH_FMIN_D            32'h2a000053
`define MASK_FMIN_D             32'hfe00707f
`define MATCH_FMAX_D            32'h2a001053
`define MASK_FMAX_D             32'hfe00707f
`define MATCH_FCVT_S_D          32'h40100053
`define MASK_FCVT_S_D           32'hfff0007f
`define MATCH_FCVT_D_S          32'h42000053
`define MASK_FCVT_D_S           32'hfff0007f
`define MATCH_FSQRT_D           32'h5a000053
`define MASK_FSQRT_D            32'hfff0007f
`define MATCH_FADD_Q            32'h6000053
`define MASK_FADD_Q             32'hfe00007f
`define MATCH_FSUB_Q            32'he000053
`define MASK_FSUB_Q             32'hfe00007f
`define MATCH_FMUL_Q            32'h16000053
`define MASK_FMUL_Q             32'hfe00007f
`define MATCH_FDIV_Q            32'h1e000053
`define MASK_FDIV_Q             32'hfe00007f
`define MATCH_FSGNJ_Q           32'h26000053
`define MASK_FSGNJ_Q            32'hfe00707f
`define MATCH_FSGNJN_Q          32'h26001053
`define MASK_FSGNJN_Q           32'hfe00707f
`define MATCH_FSGNJX_Q          32'h26002053
`define MASK_FSGNJX_Q           32'hfe00707f
`define MATCH_FMIN_Q            32'h2e000053
`define MASK_FMIN_Q             32'hfe00707f
`define MATCH_FMAX_Q            32'h2e001053
`define MASK_FMAX_Q             32'hfe00707f
`define MATCH_FCVT_S_Q          32'h40300053
`define MASK_FCVT_S_Q           32'hfff0007f
`define MATCH_FCVT_Q_S          32'h46000053
`define MASK_FCVT_Q_S           32'hfff0007f
`define MATCH_FCVT_D_Q          32'h42300053
`define MASK_FCVT_D_Q           32'hfff0007f
`define MATCH_FCVT_Q_D          32'h46100053
`define MASK_FCVT_Q_D           32'hfff0007f
`define MATCH_FSQRT_Q           32'h5e000053
`define MASK_FSQRT_Q            32'hfff0007f
`define MATCH_FLE_S             32'ha0000053
`define MASK_FLE_S              32'hfe00707f
`define MATCH_FLT_S             32'ha0001053
`define MASK_FLT_S              32'hfe00707f
`define MATCH_FEQ_S             32'ha0002053
`define MASK_FEQ_S              32'hfe00707f
`define MATCH_FLE_D             32'ha2000053
`define MASK_FLE_D              32'hfe00707f
`define MATCH_FLT_D             32'ha2001053
`define MASK_FLT_D              32'hfe00707f
`define MATCH_FEQ_D             32'ha2002053
`define MASK_FEQ_D              32'hfe00707f
`define MATCH_FLE_Q             32'ha6000053
`define MASK_FLE_Q              32'hfe00707f
`define MATCH_FLT_Q             32'ha6001053
`define MASK_FLT_Q              32'hfe00707f
`define MATCH_FEQ_Q             32'ha6002053
`define MASK_FEQ_Q              32'hfe00707f
`define MATCH_FCVT_W_S          32'hc0000053
`define MASK_FCVT_W_S           32'hfff0007f
`define MATCH_FCVT_WU_S         32'hc0100053
`define MASK_FCVT_WU_S          32'hfff0007f
`define MATCH_FCVT_L_S          32'hc0200053
`define MASK_FCVT_L_S           32'hfff0007f
`define MATCH_FCVT_LU_S         32'hc0300053
`define MASK_FCVT_LU_S          32'hfff0007f
`define MATCH_FMV_X_S           32'he0000053
`define MASK_FMV_X_S            32'hfff0707f
`define MATCH_FCLASS_S          32'he0001053
`define MASK_FCLASS_S           32'hfff0707f
`define MATCH_FCVT_W_D          32'hc2000053
`define MASK_FCVT_W_D           32'hfff0007f
`define MATCH_FCVT_WU_D         32'hc2100053
`define MASK_FCVT_WU_D          32'hfff0007f
`define MATCH_FCVT_L_D          32'hc2200053
`define MASK_FCVT_L_D           32'hfff0007f
`define MATCH_FCVT_LU_D         32'hc2300053
`define MASK_FCVT_LU_D          32'hfff0007f
`define MATCH_FMV_X_D           32'he2000053
`define MASK_FMV_X_D            32'hfff0707f
`define MATCH_FCLASS_D          32'he2001053
`define MASK_FCLASS_D           32'hfff0707f
`define MATCH_FCVT_W_Q          32'hc6000053
`define MASK_FCVT_W_Q           32'hfff0007f
`define MATCH_FCVT_WU_Q         32'hc6100053
`define MASK_FCVT_WU_Q          32'hfff0007f
`define MATCH_FCVT_L_Q          32'hc6200053
`define MASK_FCVT_L_Q           32'hfff0007f
`define MATCH_FCVT_LU_Q         32'hc6300053
`define MASK_FCVT_LU_Q          32'hfff0007f
`define MATCH_FMV_X_Q           32'he6000053
`define MASK_FMV_X_Q            32'hfff0707f
`define MATCH_FCLASS_Q          32'he6001053
`define MASK_FCLASS_Q           32'hfff0707f
`define MATCH_FCVT_S_W          32'hd0000053
`define MASK_FCVT_S_W           32'hfff0007f
`define MATCH_FCVT_S_WU         32'hd0100053
`define MASK_FCVT_S_WU          32'hfff0007f
`define MATCH_FCVT_S_L          32'hd0200053
`define MASK_FCVT_S_L           32'hfff0007f
`define MATCH_FCVT_S_LU         32'hd0300053
`define MASK_FCVT_S_LU          32'hfff0007f
`define MATCH_FMV_S_X           32'hf0000053
`define MASK_FMV_S_X            32'hfff0707f
`define MATCH_FCVT_D_W          32'hd2000053
`define MASK_FCVT_D_W           32'hfff0007f
`define MATCH_FCVT_D_WU         32'hd2100053
`define MASK_FCVT_D_WU          32'hfff0007f
`define MATCH_FCVT_D_L          32'hd2200053
`define MASK_FCVT_D_L           32'hfff0007f
`define MATCH_FCVT_D_LU         32'hd2300053
`define MASK_FCVT_D_LU          32'hfff0007f
`define MATCH_FMV_D_X           32'hf2000053
`define MASK_FMV_D_X            32'hfff0707f
`define MATCH_FCVT_Q_W          32'hd6000053
`define MASK_FCVT_Q_W           32'hfff0007f
`define MATCH_FCVT_Q_WU         32'hd6100053
`define MASK_FCVT_Q_WU          32'hfff0007f
`define MATCH_FCVT_Q_L          32'hd6200053
`define MASK_FCVT_Q_L           32'hfff0007f
`define MATCH_FCVT_Q_LU         32'hd6300053
`define MASK_FCVT_Q_LU          32'hfff0007f
`define MATCH_FMV_Q_X           32'hf6000053
`define MASK_FMV_Q_X            32'hfff0707f
`define MATCH_CLZ               32'h60001013
`define MASK_CLZ                32'hfff0707f
`define MATCH_CTZ               32'h60101013
`define MASK_CTZ                32'hfff0707f
`define MATCH_CPOP              32'h60201013
`define MASK_CPOP               32'hfff0707f
`define MATCH_MIN               32'ha004033
`define MASK_MIN                32'hfe00707f
`define MATCH_MINU              32'ha005033
`define MASK_MINU               32'hfe00707f
`define MATCH_MAX               32'ha006033
`define MASK_MAX                32'hfe00707f
`define MATCH_MAXU              32'ha007033
`define MASK_MAXU               32'hfe00707f
`define MATCH_SEXT_B            32'h60401013
`define MASK_SEXT_B             32'hfff0707f
`define MATCH_SEXT_H            32'h60501013
`define MASK_SEXT_H             32'hfff0707f
`define MATCH_PACK              32'h8004033
`define MASK_PACK               32'hfe00707f
`define MATCH_PACKH             32'h8007033
`define MASK_PACKH              32'hfe00707f
`define MATCH_PACKW             32'h800403b
`define MASK_PACKW              32'hfe00707f
`define MATCH_ANDN              32'h40007033
`define MASK_ANDN               32'hfe00707f
`define MATCH_ORN               32'h40006033
`define MASK_ORN                32'hfe00707f
`define MATCH_XNOR              32'h40004033
`define MASK_XNOR               32'hfe00707f
`define MATCH_ROL               32'h60001033
`define MASK_ROL                32'hfe00707f
`define MATCH_ROR               32'h60005033
`define MASK_ROR                32'hfe00707f
`define MATCH_RORI              32'h60005013
`define MASK_RORI               32'hfc00707f
`define MATCH_GREVI             32'h68005013
`define MASK_GREVI              32'hfc00707f
`define MATCH_GORCI             32'h28005013
`define MASK_GORCI              32'hfc00707f
`define MATCH_SHFLI             32'h8001013
`define MASK_SHFLI              32'hfe00707f
`define MATCH_UNSHFLI           32'h8005013
`define MASK_UNSHFLI            32'hfe00707f
`define MATCH_CLZW              32'h6000101b
`define MASK_CLZW               32'hfff0707f
`define MATCH_CTZW              32'h6010101b
`define MASK_CTZW               32'hfff0707f
`define MATCH_CPOPW             32'h6020101b
`define MASK_CPOPW              32'hfff0707f
`define MATCH_ROLW              32'h6000103b
`define MASK_ROLW               32'hfe00707f
`define MATCH_RORW              32'h6000503b
`define MASK_RORW               32'hfe00707f
`define MATCH_RORIW             32'h6000501b
`define MASK_RORIW              32'hfe00707f
`define MATCH_SH1ADD            32'h20002033
`define MASK_SH1ADD             32'hfe00707f
`define MATCH_SH2ADD            32'h20004033
`define MASK_SH2ADD             32'hfe00707f
`define MATCH_SH3ADD            32'h20006033
`define MASK_SH3ADD             32'hfe00707f
`define MATCH_SH1ADD_UW         32'h2000203b
`define MASK_SH1ADD_UW          32'hfe00707f
`define MATCH_SH2ADD_UW         32'h2000403b
`define MASK_SH2ADD_UW          32'hfe00707f
`define MATCH_SH3ADD_UW         32'h2000603b
`define MASK_SH3ADD_UW          32'hfe00707f
`define MATCH_ADD_UW            32'h800003b
`define MASK_ADD_UW             32'hfe00707f
`define MATCH_SLLI_UW           32'h800101b
`define MASK_SLLI_UW            32'hfc00707f
`define MATCH_CLMUL             32'ha001033
`define MASK_CLMUL              32'hfe00707f
`define MATCH_CLMULH            32'ha003033
`define MASK_CLMULH             32'hfe00707f
`define MATCH_CLMULR            32'ha002033
`define MASK_CLMULR             32'hfe00707f
`define MATCH_XPERM4            32'h28002033
`define MASK_XPERM4             32'hfe00707f
`define MATCH_XPERM8            32'h28004033
`define MASK_XPERM8             32'hfe00707f
`define MATCH_BCLRI             32'h48001013
`define MASK_BCLRI              32'hfc00707f
`define MATCH_BSETI             32'h28001013
`define MASK_BSETI              32'hfc00707f
`define MATCH_BINVI             32'h68001013
`define MASK_BINVI              32'hfc00707f
`define MATCH_BEXTI             32'h48005013
`define MASK_BEXTI              32'hfc00707f
`define MATCH_BCLR              32'h48001033
`define MASK_BCLR               32'hfe00707f
`define MATCH_BSET              32'h28001033
`define MASK_BSET               32'hfe00707f
`define MATCH_BINV              32'h68001033
`define MASK_BINV               32'hfe00707f
`define MATCH_BEXT              32'h48005033
`define MASK_BEXT               32'hfe00707f
`define MATCH_FLW               32'h2007
`define MASK_FLW                32'h707f
`define MATCH_FLD               32'h3007
`define MASK_FLD                32'h707f
`define MATCH_FLQ               32'h4007
`define MASK_FLQ                32'h707f
`define MATCH_FSW               32'h2027
`define MASK_FSW                32'h707f
`define MATCH_FSD               32'h3027
`define MASK_FSD                32'h707f
`define MATCH_FSQ               32'h4027
`define MASK_FSQ                32'h707f
`define MATCH_FMADD_S           32'h43
`define MASK_FMADD_S            32'h600007f
`define MATCH_FMSUB_S           32'h47
`define MASK_FMSUB_S            32'h600007f
`define MATCH_FNMSUB_S          32'h4b
`define MASK_FNMSUB_S           32'h600007f
`define MATCH_FNMADD_S          32'h4f
`define MASK_FNMADD_S           32'h600007f
`define MATCH_FMADD_D           32'h2000043
`define MASK_FMADD_D            32'h600007f
`define MATCH_FMSUB_D           32'h2000047
`define MASK_FMSUB_D            32'h600007f
`define MATCH_FNMSUB_D          32'h200004b
`define MASK_FNMSUB_D           32'h600007f
`define MATCH_FNMADD_D          32'h200004f
`define MASK_FNMADD_D           32'h600007f
`define MATCH_FMADD_Q           32'h6000043
`define MASK_FMADD_Q            32'h600007f
`define MATCH_FMSUB_Q           32'h6000047
`define MASK_FMSUB_Q            32'h600007f
`define MATCH_FNMSUB_Q          32'h600004b
`define MASK_FNMSUB_Q           32'h600007f
`define MATCH_FNMADD_Q          32'h600004f
`define MASK_FNMADD_Q           32'h600007f
`define MATCH_C_ADDI4SPN        32'h0
`define MASK_C_ADDI4SPN         32'he003
`define MATCH_C_FLD             32'h2000
`define MASK_C_FLD              32'he003
`define MATCH_C_LW              32'h4000
`define MASK_C_LW               32'he003
`define MATCH_C_FLW             32'h6000
`define MASK_C_FLW              32'he003
`define MATCH_C_FSD             32'ha000
`define MASK_C_FSD              32'he003
`define MATCH_C_SW              32'hc000
`define MASK_C_SW               32'he003
`define MATCH_C_FSW             32'he000
`define MASK_C_FSW              32'he003
`define MATCH_C_ADDI            32'h1
`define MASK_C_ADDI             32'he003
`define MATCH_C_JAL             32'h2001
`define MASK_C_JAL              32'he003
`define MATCH_C_LI              32'h4001
`define MASK_C_LI               32'he003
`define MATCH_C_LUI             32'h6001
`define MASK_C_LUI              32'he003
`define MATCH_C_SRLI            32'h8001
`define MASK_C_SRLI             32'hec03
`define MATCH_C_SRLI64          32'h8001
`define MASK_C_SRLI64           32'hfc7f
`define MATCH_C_SRAI            32'h8401
`define MASK_C_SRAI             32'hec03
`define MATCH_C_SRAI64          32'h8401
`define MASK_C_SRAI64           32'hfc7f
`define MATCH_C_ANDI            32'h8801
`define MASK_C_ANDI             32'hec03
`define MATCH_C_SUB             32'h8c01
`define MASK_C_SUB              32'hfc63
`define MATCH_C_XOR             32'h8c21
`define MASK_C_XOR              32'hfc63
`define MATCH_C_OR              32'h8c41
`define MASK_C_OR               32'hfc63
`define MATCH_C_AND             32'h8c61
`define MASK_C_AND              32'hfc63
`define MATCH_C_SUBW            32'h9c01
`define MASK_C_SUBW             32'hfc63
`define MATCH_C_ADDW            32'h9c21
`define MASK_C_ADDW             32'hfc63
`define MATCH_C_J               32'ha001
`define MASK_C_J                32'he003
`define MATCH_C_BEQZ            32'hc001
`define MASK_C_BEQZ             32'he003
`define MATCH_C_BNEZ            32'he001
`define MASK_C_BNEZ             32'he003
`define MATCH_C_SLLI            32'h2
`define MASK_C_SLLI             32'he003
`define MATCH_C_SLLI64          32'h2
`define MASK_C_SLLI64           32'hf07f
`define MATCH_C_FLDSP           32'h2002
`define MASK_C_FLDSP            32'he003
`define MATCH_C_LWSP            32'h4002
`define MASK_C_LWSP             32'he003
`define MATCH_C_FLWSP           32'h6002
`define MASK_C_FLWSP            32'he003
`define MATCH_C_MV              32'h8002
`define MASK_C_MV               32'hf003
`define MATCH_C_ADD             32'h9002
`define MASK_C_ADD              32'hf003
`define MATCH_C_FSDSP           32'ha002
`define MASK_C_FSDSP            32'he003
`define MATCH_C_SWSP            32'hc002
`define MASK_C_SWSP             32'he003
`define MATCH_C_FSWSP           32'he002
`define MASK_C_FSWSP            32'he003
`define MATCH_C_NOP             32'h1
`define MASK_C_NOP              32'hffff
`define MATCH_C_ADDI16SP        32'h6101
`define MASK_C_ADDI16SP         32'hef83
`define MATCH_C_JR              32'h8002
`define MASK_C_JR               32'hf07f
`define MATCH_C_JALR            32'h9002
`define MASK_C_JALR             32'hf07f
`define MATCH_C_EBREAK          32'h9002
`define MASK_C_EBREAK           32'hffff
`define MATCH_C_LD              32'h6000
`define MASK_C_LD               32'he003
`define MATCH_C_SD              32'he000
`define MASK_C_SD               32'he003
`define MATCH_C_ADDIW           32'h2001
`define MASK_C_ADDIW            32'he003
`define MATCH_C_LDSP            32'h6002
`define MASK_C_LDSP             32'he003
`define MATCH_C_SDSP            32'he002
`define MASK_C_SDSP             32'he003