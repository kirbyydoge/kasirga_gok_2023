`timescale 1ns/1ps

`include "sabitler.vh"
`include "mikroislem.vh"

module veri_yolu_birimi(
    input                      clk_i,
    input                      rstn_i,

    input   [`UOP_BEL_BIT-1:0] uop_buyruk_secim_i,
    input   [`UOP_RS1_BIT-1:0] uop_rs1_i,
    input   [`UOP_RS2_BIT-1:0] uop_rs2_i,
    input   [`UOP_IMM_BIT-1:0] uop_imm_i

    //YAZILACAK (ŞEVVAL) 

       
);
endmodule